module digel_soc (clk,
    flash_clk,
    flash_csb,
    flash_io0,
    flash_io1,
    flash_io2,
    flash_io3,
    led1,
    led2,
    led3,
    led4,
    led5,
    ledg_n,
    ledr_n,
    ser_rx,
    ser_tx,
    mode,
    wave);
 input clk;
 output flash_clk;
 output flash_csb;
 inout flash_io0;
 inout flash_io1;
 inout flash_io2;
 inout flash_io3;
 output led1;
 output led2;
 output led3;
 output led4;
 output led5;
 output ledg_n;
 output ledr_n;
 input ser_rx;
 output ser_tx;
 output [2:0] mode;
 output [31:0] wave;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _146_;
 wire _147_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire net419;
 wire flash_io0_oe;
 wire flash_io1_oe;
 wire flash_io2_oe;
 wire flash_io3_oe;
 wire \gpio[0] ;
 wire \gpio[10] ;
 wire \gpio[11] ;
 wire \gpio[12] ;
 wire \gpio[13] ;
 wire \gpio[14] ;
 wire \gpio[15] ;
 wire \gpio[16] ;
 wire \gpio[17] ;
 wire \gpio[18] ;
 wire \gpio[19] ;
 wire \gpio[20] ;
 wire \gpio[21] ;
 wire \gpio[22] ;
 wire \gpio[23] ;
 wire \gpio[24] ;
 wire \gpio[25] ;
 wire \gpio[26] ;
 wire \gpio[27] ;
 wire \gpio[28] ;
 wire \gpio[29] ;
 wire \gpio[30] ;
 wire \gpio[31] ;
 wire \gpio[6] ;
 wire \gpio[7] ;
 wire \gpio[8] ;
 wire \gpio[9] ;
 wire net712;
 wire \iomem_addr[10] ;
 wire \iomem_addr[11] ;
 wire \iomem_addr[12] ;
 wire \iomem_addr[13] ;
 wire \iomem_addr[14] ;
 wire \iomem_addr[15] ;
 wire \iomem_addr[16] ;
 wire \iomem_addr[17] ;
 wire \iomem_addr[18] ;
 wire \iomem_addr[19] ;
 wire net711;
 wire \iomem_addr[20] ;
 wire \iomem_addr[21] ;
 wire \iomem_addr[22] ;
 wire \iomem_addr[23] ;
 wire \iomem_addr[24] ;
 wire \iomem_addr[25] ;
 wire \iomem_addr[26] ;
 wire \iomem_addr[27] ;
 wire \iomem_addr[28] ;
 wire \iomem_addr[29] ;
 wire \iomem_addr[2] ;
 wire \iomem_addr[30] ;
 wire \iomem_addr[31] ;
 wire \iomem_addr[3] ;
 wire \iomem_addr[4] ;
 wire \iomem_addr[5] ;
 wire \iomem_addr[6] ;
 wire \iomem_addr[7] ;
 wire \iomem_addr[8] ;
 wire \iomem_addr[9] ;
 wire \iomem_rdata[0] ;
 wire \iomem_rdata[10] ;
 wire \iomem_rdata[11] ;
 wire \iomem_rdata[12] ;
 wire \iomem_rdata[13] ;
 wire \iomem_rdata[14] ;
 wire \iomem_rdata[15] ;
 wire \iomem_rdata[16] ;
 wire \iomem_rdata[17] ;
 wire \iomem_rdata[18] ;
 wire \iomem_rdata[19] ;
 wire \iomem_rdata[1] ;
 wire \iomem_rdata[20] ;
 wire \iomem_rdata[21] ;
 wire \iomem_rdata[22] ;
 wire \iomem_rdata[23] ;
 wire \iomem_rdata[24] ;
 wire \iomem_rdata[25] ;
 wire \iomem_rdata[26] ;
 wire \iomem_rdata[27] ;
 wire \iomem_rdata[28] ;
 wire \iomem_rdata[29] ;
 wire \iomem_rdata[2] ;
 wire \iomem_rdata[30] ;
 wire \iomem_rdata[31] ;
 wire \iomem_rdata[3] ;
 wire \iomem_rdata[4] ;
 wire \iomem_rdata[5] ;
 wire \iomem_rdata[6] ;
 wire \iomem_rdata[7] ;
 wire \iomem_rdata[8] ;
 wire \iomem_rdata[9] ;
 wire iomem_ready;
 wire iomem_valid;
 wire \iomem_wdata[0] ;
 wire \iomem_wdata[10] ;
 wire \iomem_wdata[11] ;
 wire \iomem_wdata[12] ;
 wire \iomem_wdata[13] ;
 wire \iomem_wdata[14] ;
 wire \iomem_wdata[15] ;
 wire \iomem_wdata[16] ;
 wire \iomem_wdata[17] ;
 wire \iomem_wdata[18] ;
 wire \iomem_wdata[19] ;
 wire \iomem_wdata[1] ;
 wire \iomem_wdata[20] ;
 wire \iomem_wdata[21] ;
 wire \iomem_wdata[22] ;
 wire \iomem_wdata[23] ;
 wire \iomem_wdata[24] ;
 wire \iomem_wdata[25] ;
 wire \iomem_wdata[26] ;
 wire \iomem_wdata[27] ;
 wire \iomem_wdata[28] ;
 wire \iomem_wdata[29] ;
 wire \iomem_wdata[2] ;
 wire \iomem_wdata[30] ;
 wire \iomem_wdata[31] ;
 wire \iomem_wdata[3] ;
 wire \iomem_wdata[4] ;
 wire \iomem_wdata[5] ;
 wire \iomem_wdata[6] ;
 wire \iomem_wdata[7] ;
 wire \iomem_wdata[8] ;
 wire \iomem_wdata[9] ;
 wire \iomem_wstrb[0] ;
 wire \iomem_wstrb[1] ;
 wire \iomem_wstrb[2] ;
 wire \iomem_wstrb[3] ;
 wire \reset_cnt[0] ;
 wire \reset_cnt[1] ;
 wire \reset_cnt[2] ;
 wire \reset_cnt[3] ;
 wire \reset_cnt[4] ;
 wire \reset_cnt[5] ;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire \soc/_000_ ;
 wire \soc/_001_ ;
 wire \soc/_002_ ;
 wire \soc/_003_ ;
 wire \soc/_004_ ;
 wire \soc/_005_ ;
 wire \soc/_006_ ;
 wire \soc/_007_ ;
 wire \soc/_008_ ;
 wire \soc/_009_ ;
 wire \soc/_010_ ;
 wire \soc/_011_ ;
 wire \soc/_012_ ;
 wire \soc/_013_ ;
 wire \soc/_014_ ;
 wire \soc/_015_ ;
 wire \soc/_016_ ;
 wire \soc/_017_ ;
 wire \soc/_018_ ;
 wire \soc/_019_ ;
 wire \soc/_020_ ;
 wire \soc/_021_ ;
 wire \soc/_022_ ;
 wire \soc/_023_ ;
 wire \soc/_024_ ;
 wire \soc/_025_ ;
 wire \soc/_026_ ;
 wire \soc/_027_ ;
 wire \soc/_028_ ;
 wire \soc/_029_ ;
 wire \soc/_030_ ;
 wire \soc/_031_ ;
 wire \soc/_032_ ;
 wire \soc/_033_ ;
 wire \soc/_034_ ;
 wire \soc/_036_ ;
 wire \soc/_037_ ;
 wire \soc/_039_ ;
 wire \soc/_040_ ;
 wire \soc/_041_ ;
 wire \soc/_042_ ;
 wire \soc/_044_ ;
 wire \soc/_049_ ;
 wire \soc/_053_ ;
 wire \soc/_054_ ;
 wire \soc/_056_ ;
 wire \soc/_058_ ;
 wire \soc/_059_ ;
 wire \soc/_060_ ;
 wire \soc/_061_ ;
 wire \soc/_062_ ;
 wire \soc/_063_ ;
 wire \soc/_064_ ;
 wire \soc/_065_ ;
 wire \soc/_066_ ;
 wire \soc/_067_ ;
 wire \soc/_068_ ;
 wire \soc/_069_ ;
 wire \soc/_070_ ;
 wire \soc/_071_ ;
 wire \soc/_072_ ;
 wire \soc/_073_ ;
 wire \soc/_074_ ;
 wire \soc/_075_ ;
 wire \soc/_076_ ;
 wire \soc/_077_ ;
 wire \soc/_078_ ;
 wire \soc/_081_ ;
 wire \soc/_082_ ;
 wire \soc/_083_ ;
 wire \soc/_084_ ;
 wire \soc/_085_ ;
 wire \soc/_086_ ;
 wire \soc/_087_ ;
 wire \soc/_088_ ;
 wire \soc/_089_ ;
 wire \soc/_090_ ;
 wire \soc/_091_ ;
 wire \soc/_092_ ;
 wire \soc/_093_ ;
 wire \soc/_094_ ;
 wire \soc/_095_ ;
 wire \soc/_097_ ;
 wire \soc/_100_ ;
 wire \soc/_101_ ;
 wire \soc/_102_ ;
 wire \soc/_104_ ;
 wire \soc/_105_ ;
 wire \soc/_106_ ;
 wire \soc/_107_ ;
 wire \soc/_108_ ;
 wire \soc/_109_ ;
 wire \soc/_112_ ;
 wire \soc/_113_ ;
 wire \soc/_114_ ;
 wire \soc/_116_ ;
 wire \soc/_117_ ;
 wire \soc/_118_ ;
 wire \soc/_119_ ;
 wire \soc/_120_ ;
 wire \soc/_121_ ;
 wire \soc/_122_ ;
 wire \soc/_123_ ;
 wire \soc/_124_ ;
 wire \soc/_125_ ;
 wire \soc/_126_ ;
 wire \soc/_127_ ;
 wire \soc/_128_ ;
 wire \soc/_129_ ;
 wire \soc/_130_ ;
 wire \soc/_131_ ;
 wire \soc/_132_ ;
 wire \soc/_133_ ;
 wire \soc/_134_ ;
 wire \soc/_135_ ;
 wire \soc/_136_ ;
 wire \soc/_137_ ;
 wire \soc/_140_ ;
 wire \soc/_141_ ;
 wire \soc/_142_ ;
 wire \soc/_143_ ;
 wire \soc/_144_ ;
 wire \soc/_145_ ;
 wire \soc/_146_ ;
 wire \soc/_147_ ;
 wire \soc/_148_ ;
 wire \soc/_149_ ;
 wire \soc/_150_ ;
 wire \soc/_151_ ;
 wire \soc/_152_ ;
 wire \soc/_153_ ;
 wire \soc/_154_ ;
 wire \soc/_156_ ;
 wire \soc/_159_ ;
 wire \soc/_160_ ;
 wire \soc/_161_ ;
 wire \soc/_163_ ;
 wire \soc/_164_ ;
 wire \soc/_165_ ;
 wire \soc/_166_ ;
 wire \soc/_167_ ;
 wire \soc/_168_ ;
 wire \soc/_171_ ;
 wire \soc/_172_ ;
 wire \soc/_173_ ;
 wire \soc/_175_ ;
 wire \soc/_176_ ;
 wire \soc/_177_ ;
 wire \soc/_178_ ;
 wire \soc/_179_ ;
 wire \soc/_180_ ;
 wire \soc/_181_ ;
 wire \soc/_182_ ;
 wire \soc/_183_ ;
 wire \soc/_184_ ;
 wire \soc/_185_ ;
 wire \soc/_186_ ;
 wire \soc/_187_ ;
 wire \soc/_188_ ;
 wire \soc/_189_ ;
 wire \soc/_190_ ;
 wire \soc/_191_ ;
 wire \soc/_192_ ;
 wire \soc/_193_ ;
 wire \soc/_194_ ;
 wire \soc/_195_ ;
 wire \soc/_196_ ;
 wire \soc/_197_ ;
 wire \soc/_198_ ;
 wire \soc/_199_ ;
 wire \soc/_200_ ;
 wire \soc/_201_ ;
 wire \soc/_202_ ;
 wire \soc/_203_ ;
 wire \soc/_204_ ;
 wire \soc/_205_ ;
 wire \soc/_206_ ;
 wire \soc/_207_ ;
 wire \soc/_208_ ;
 wire \soc/_209_ ;
 wire \soc/_210_ ;
 wire \soc/_211_ ;
 wire \soc/_212_ ;
 wire \soc/_213_ ;
 wire \soc/_214_ ;
 wire \soc/_215_ ;
 wire \soc/_216_ ;
 wire \soc/_217_ ;
 wire \soc/_218_ ;
 wire \soc/_219_ ;
 wire \soc/_220_ ;
 wire \soc/_221_ ;
 wire \soc/_222_ ;
 wire \soc/_223_ ;
 wire \soc/_224_ ;
 wire \soc/_225_ ;
 wire \soc/_226_ ;
 wire \soc/_227_ ;
 wire \soc/_228_ ;
 wire \soc/_229_ ;
 wire \soc/_230_ ;
 wire \soc/_231_ ;
 wire net448;
 wire \soc/mem_instr ;
 wire \soc/mem_rdata[0] ;
 wire \soc/mem_rdata[10] ;
 wire \soc/mem_rdata[11] ;
 wire \soc/mem_rdata[12] ;
 wire \soc/mem_rdata[13] ;
 wire \soc/mem_rdata[14] ;
 wire \soc/mem_rdata[15] ;
 wire \soc/mem_rdata[16] ;
 wire \soc/mem_rdata[17] ;
 wire \soc/mem_rdata[18] ;
 wire \soc/mem_rdata[19] ;
 wire \soc/mem_rdata[1] ;
 wire \soc/mem_rdata[20] ;
 wire \soc/mem_rdata[21] ;
 wire \soc/mem_rdata[22] ;
 wire \soc/mem_rdata[23] ;
 wire \soc/mem_rdata[24] ;
 wire \soc/mem_rdata[25] ;
 wire \soc/mem_rdata[26] ;
 wire \soc/mem_rdata[27] ;
 wire \soc/mem_rdata[28] ;
 wire \soc/mem_rdata[29] ;
 wire \soc/mem_rdata[2] ;
 wire \soc/mem_rdata[30] ;
 wire \soc/mem_rdata[31] ;
 wire \soc/mem_rdata[3] ;
 wire \soc/mem_rdata[4] ;
 wire \soc/mem_rdata[5] ;
 wire \soc/mem_rdata[6] ;
 wire \soc/mem_rdata[7] ;
 wire \soc/mem_rdata[8] ;
 wire \soc/mem_rdata[9] ;
 wire \soc/mem_ready ;
 wire \soc/mem_valid ;
 wire \soc/ram_rdata[0] ;
 wire \soc/ram_rdata[10] ;
 wire \soc/ram_rdata[11] ;
 wire \soc/ram_rdata[12] ;
 wire \soc/ram_rdata[13] ;
 wire \soc/ram_rdata[14] ;
 wire \soc/ram_rdata[15] ;
 wire \soc/ram_rdata[16] ;
 wire \soc/ram_rdata[17] ;
 wire \soc/ram_rdata[18] ;
 wire \soc/ram_rdata[19] ;
 wire \soc/ram_rdata[1] ;
 wire \soc/ram_rdata[20] ;
 wire \soc/ram_rdata[21] ;
 wire \soc/ram_rdata[22] ;
 wire \soc/ram_rdata[23] ;
 wire \soc/ram_rdata[24] ;
 wire \soc/ram_rdata[25] ;
 wire \soc/ram_rdata[26] ;
 wire \soc/ram_rdata[27] ;
 wire \soc/ram_rdata[28] ;
 wire \soc/ram_rdata[29] ;
 wire \soc/ram_rdata[2] ;
 wire \soc/ram_rdata[30] ;
 wire \soc/ram_rdata[31] ;
 wire \soc/ram_rdata[3] ;
 wire \soc/ram_rdata[4] ;
 wire \soc/ram_rdata[5] ;
 wire \soc/ram_rdata[6] ;
 wire \soc/ram_rdata[7] ;
 wire \soc/ram_rdata[8] ;
 wire \soc/ram_rdata[9] ;
 wire \soc/ram_ready ;
 wire \soc/simpleuart_reg_dat_do[0] ;
 wire net320;
 wire net319;
 wire net318;
 wire net317;
 wire net316;
 wire net315;
 wire net314;
 wire net313;
 wire net312;
 wire net311;
 wire \soc/simpleuart_reg_dat_do[1] ;
 wire net310;
 wire net309;
 wire net308;
 wire net307;
 wire net306;
 wire net305;
 wire net304;
 wire net303;
 wire net302;
 wire net301;
 wire \soc/simpleuart_reg_dat_do[2] ;
 wire net300;
 wire \soc/simpleuart_reg_dat_do[31] ;
 wire \soc/simpleuart_reg_dat_do[3] ;
 wire \soc/simpleuart_reg_dat_do[4] ;
 wire \soc/simpleuart_reg_dat_do[5] ;
 wire \soc/simpleuart_reg_dat_do[6] ;
 wire \soc/simpleuart_reg_dat_do[7] ;
 wire net322;
 wire net321;
 wire \soc/simpleuart_reg_dat_wait ;
 wire \soc/simpleuart_reg_div_do[0] ;
 wire \soc/simpleuart_reg_div_do[10] ;
 wire \soc/simpleuart_reg_div_do[11] ;
 wire \soc/simpleuart_reg_div_do[12] ;
 wire \soc/simpleuart_reg_div_do[13] ;
 wire \soc/simpleuart_reg_div_do[14] ;
 wire \soc/simpleuart_reg_div_do[15] ;
 wire \soc/simpleuart_reg_div_do[16] ;
 wire \soc/simpleuart_reg_div_do[17] ;
 wire \soc/simpleuart_reg_div_do[18] ;
 wire \soc/simpleuart_reg_div_do[19] ;
 wire \soc/simpleuart_reg_div_do[1] ;
 wire \soc/simpleuart_reg_div_do[20] ;
 wire \soc/simpleuart_reg_div_do[21] ;
 wire \soc/simpleuart_reg_div_do[22] ;
 wire \soc/simpleuart_reg_div_do[23] ;
 wire \soc/simpleuart_reg_div_do[24] ;
 wire \soc/simpleuart_reg_div_do[25] ;
 wire \soc/simpleuart_reg_div_do[26] ;
 wire \soc/simpleuart_reg_div_do[27] ;
 wire \soc/simpleuart_reg_div_do[28] ;
 wire \soc/simpleuart_reg_div_do[29] ;
 wire \soc/simpleuart_reg_div_do[2] ;
 wire \soc/simpleuart_reg_div_do[30] ;
 wire \soc/simpleuart_reg_div_do[31] ;
 wire \soc/simpleuart_reg_div_do[3] ;
 wire \soc/simpleuart_reg_div_do[4] ;
 wire \soc/simpleuart_reg_div_do[5] ;
 wire \soc/simpleuart_reg_div_do[6] ;
 wire \soc/simpleuart_reg_div_do[7] ;
 wire \soc/simpleuart_reg_div_do[8] ;
 wire \soc/simpleuart_reg_div_do[9] ;
 wire \soc/spimem_rdata[0] ;
 wire \soc/spimem_rdata[10] ;
 wire \soc/spimem_rdata[11] ;
 wire \soc/spimem_rdata[12] ;
 wire \soc/spimem_rdata[13] ;
 wire \soc/spimem_rdata[14] ;
 wire \soc/spimem_rdata[15] ;
 wire \soc/spimem_rdata[16] ;
 wire \soc/spimem_rdata[17] ;
 wire \soc/spimem_rdata[18] ;
 wire \soc/spimem_rdata[19] ;
 wire \soc/spimem_rdata[1] ;
 wire \soc/spimem_rdata[20] ;
 wire \soc/spimem_rdata[21] ;
 wire \soc/spimem_rdata[22] ;
 wire \soc/spimem_rdata[23] ;
 wire \soc/spimem_rdata[24] ;
 wire \soc/spimem_rdata[25] ;
 wire \soc/spimem_rdata[26] ;
 wire \soc/spimem_rdata[27] ;
 wire \soc/spimem_rdata[28] ;
 wire \soc/spimem_rdata[29] ;
 wire \soc/spimem_rdata[2] ;
 wire \soc/spimem_rdata[30] ;
 wire \soc/spimem_rdata[31] ;
 wire \soc/spimem_rdata[3] ;
 wire \soc/spimem_rdata[4] ;
 wire \soc/spimem_rdata[5] ;
 wire \soc/spimem_rdata[6] ;
 wire \soc/spimem_rdata[7] ;
 wire \soc/spimem_rdata[8] ;
 wire \soc/spimem_rdata[9] ;
 wire \soc/spimem_ready ;
 wire net269;
 wire net259;
 wire net258;
 wire net257;
 wire net256;
 wire net255;
 wire net254;
 wire \soc/spimemio_cfgreg_do[16] ;
 wire \soc/spimemio_cfgreg_do[17] ;
 wire \soc/spimemio_cfgreg_do[18] ;
 wire \soc/spimemio_cfgreg_do[19] ;
 wire net268;
 wire net253;
 wire net252;
 wire net251;
 wire net250;
 wire net249;
 wire net248;
 wire net247;
 wire net246;
 wire net245;
 wire net244;
 wire net267;
 wire net243;
 wire net242;
 wire net266;
 wire net265;
 wire net264;
 wire net263;
 wire net262;
 wire net261;
 wire net260;
 wire \soc/cpu/_00000_ ;
 wire \soc/cpu/_00001_ ;
 wire \soc/cpu/_00002_ ;
 wire \soc/cpu/_00003_ ;
 wire \soc/cpu/_00004_ ;
 wire \soc/cpu/_00005_ ;
 wire \soc/cpu/_00006_ ;
 wire \soc/cpu/_00007_ ;
 wire \soc/cpu/_00008_ ;
 wire \soc/cpu/_00009_ ;
 wire \soc/cpu/_00010_ ;
 wire \soc/cpu/_00011_ ;
 wire \soc/cpu/_00012_ ;
 wire \soc/cpu/_00013_ ;
 wire \soc/cpu/_00014_ ;
 wire \soc/cpu/_00015_ ;
 wire \soc/cpu/_00016_ ;
 wire \soc/cpu/_00017_ ;
 wire \soc/cpu/_00018_ ;
 wire \soc/cpu/_00019_ ;
 wire \soc/cpu/_00020_ ;
 wire \soc/cpu/_00021_ ;
 wire \soc/cpu/_00022_ ;
 wire \soc/cpu/_00023_ ;
 wire \soc/cpu/_00024_ ;
 wire \soc/cpu/_00025_ ;
 wire \soc/cpu/_00026_ ;
 wire \soc/cpu/_00027_ ;
 wire \soc/cpu/_00028_ ;
 wire \soc/cpu/_00029_ ;
 wire \soc/cpu/_00030_ ;
 wire \soc/cpu/_00031_ ;
 wire \soc/cpu/_00032_ ;
 wire \soc/cpu/_00033_ ;
 wire \soc/cpu/_00034_ ;
 wire \soc/cpu/_00035_ ;
 wire \soc/cpu/_00036_ ;
 wire \soc/cpu/_00037_ ;
 wire \soc/cpu/_00038_ ;
 wire \soc/cpu/_00039_ ;
 wire \soc/cpu/_00040_ ;
 wire \soc/cpu/_00041_ ;
 wire \soc/cpu/_00042_ ;
 wire \soc/cpu/_00043_ ;
 wire \soc/cpu/_00044_ ;
 wire \soc/cpu/_00045_ ;
 wire \soc/cpu/_00046_ ;
 wire \soc/cpu/_00047_ ;
 wire \soc/cpu/_00048_ ;
 wire \soc/cpu/_00049_ ;
 wire \soc/cpu/_00050_ ;
 wire \soc/cpu/_00051_ ;
 wire \soc/cpu/_00052_ ;
 wire \soc/cpu/_00053_ ;
 wire \soc/cpu/_00054_ ;
 wire \soc/cpu/_00055_ ;
 wire \soc/cpu/_00056_ ;
 wire \soc/cpu/_00057_ ;
 wire \soc/cpu/_00058_ ;
 wire \soc/cpu/_00059_ ;
 wire \soc/cpu/_00060_ ;
 wire \soc/cpu/_00061_ ;
 wire \soc/cpu/_00062_ ;
 wire \soc/cpu/_00063_ ;
 wire \soc/cpu/_00064_ ;
 wire \soc/cpu/_00065_ ;
 wire \soc/cpu/_00066_ ;
 wire \soc/cpu/_00067_ ;
 wire \soc/cpu/_00068_ ;
 wire \soc/cpu/_00069_ ;
 wire \soc/cpu/_00070_ ;
 wire \soc/cpu/_00071_ ;
 wire \soc/cpu/_00072_ ;
 wire \soc/cpu/_00073_ ;
 wire \soc/cpu/_00074_ ;
 wire \soc/cpu/_00075_ ;
 wire \soc/cpu/_00076_ ;
 wire \soc/cpu/_00077_ ;
 wire \soc/cpu/_00078_ ;
 wire \soc/cpu/_00079_ ;
 wire \soc/cpu/_00080_ ;
 wire \soc/cpu/_00081_ ;
 wire \soc/cpu/_00082_ ;
 wire \soc/cpu/_00083_ ;
 wire \soc/cpu/_00084_ ;
 wire \soc/cpu/_00085_ ;
 wire \soc/cpu/_00086_ ;
 wire \soc/cpu/_00087_ ;
 wire \soc/cpu/_00088_ ;
 wire \soc/cpu/_00089_ ;
 wire \soc/cpu/_00090_ ;
 wire \soc/cpu/_00091_ ;
 wire \soc/cpu/_00092_ ;
 wire \soc/cpu/_00093_ ;
 wire \soc/cpu/_00094_ ;
 wire \soc/cpu/_00095_ ;
 wire \soc/cpu/_00096_ ;
 wire \soc/cpu/_00097_ ;
 wire \soc/cpu/_00098_ ;
 wire \soc/cpu/_00099_ ;
 wire \soc/cpu/_00100_ ;
 wire \soc/cpu/_00101_ ;
 wire \soc/cpu/_00102_ ;
 wire \soc/cpu/_00103_ ;
 wire \soc/cpu/_00104_ ;
 wire \soc/cpu/_00105_ ;
 wire \soc/cpu/_00106_ ;
 wire \soc/cpu/_00107_ ;
 wire \soc/cpu/_00108_ ;
 wire \soc/cpu/_00109_ ;
 wire \soc/cpu/_00110_ ;
 wire \soc/cpu/_00111_ ;
 wire \soc/cpu/_00112_ ;
 wire \soc/cpu/_00113_ ;
 wire \soc/cpu/_00114_ ;
 wire \soc/cpu/_00115_ ;
 wire \soc/cpu/_00116_ ;
 wire \soc/cpu/_00117_ ;
 wire \soc/cpu/_00118_ ;
 wire \soc/cpu/_00119_ ;
 wire \soc/cpu/_00120_ ;
 wire \soc/cpu/_00121_ ;
 wire \soc/cpu/_00122_ ;
 wire \soc/cpu/_00123_ ;
 wire \soc/cpu/_00124_ ;
 wire \soc/cpu/_00125_ ;
 wire \soc/cpu/_00126_ ;
 wire \soc/cpu/_00127_ ;
 wire \soc/cpu/_00128_ ;
 wire \soc/cpu/_00129_ ;
 wire \soc/cpu/_00130_ ;
 wire \soc/cpu/_00131_ ;
 wire \soc/cpu/_00132_ ;
 wire \soc/cpu/_00133_ ;
 wire \soc/cpu/_00134_ ;
 wire \soc/cpu/_00135_ ;
 wire \soc/cpu/_00136_ ;
 wire \soc/cpu/_00137_ ;
 wire \soc/cpu/_00138_ ;
 wire \soc/cpu/_00139_ ;
 wire \soc/cpu/_00140_ ;
 wire \soc/cpu/_00141_ ;
 wire \soc/cpu/_00142_ ;
 wire \soc/cpu/_00143_ ;
 wire \soc/cpu/_00144_ ;
 wire \soc/cpu/_00145_ ;
 wire \soc/cpu/_00146_ ;
 wire \soc/cpu/_00147_ ;
 wire \soc/cpu/_00148_ ;
 wire \soc/cpu/_00149_ ;
 wire \soc/cpu/_00150_ ;
 wire \soc/cpu/_00151_ ;
 wire \soc/cpu/_00152_ ;
 wire \soc/cpu/_00153_ ;
 wire \soc/cpu/_00154_ ;
 wire \soc/cpu/_00155_ ;
 wire \soc/cpu/_00156_ ;
 wire \soc/cpu/_00157_ ;
 wire \soc/cpu/_00158_ ;
 wire \soc/cpu/_00159_ ;
 wire \soc/cpu/_00160_ ;
 wire \soc/cpu/_00161_ ;
 wire \soc/cpu/_00162_ ;
 wire \soc/cpu/_00163_ ;
 wire \soc/cpu/_00164_ ;
 wire \soc/cpu/_00165_ ;
 wire \soc/cpu/_00166_ ;
 wire \soc/cpu/_00167_ ;
 wire \soc/cpu/_00168_ ;
 wire \soc/cpu/_00169_ ;
 wire \soc/cpu/_00170_ ;
 wire \soc/cpu/_00171_ ;
 wire \soc/cpu/_00172_ ;
 wire \soc/cpu/_00173_ ;
 wire \soc/cpu/_00174_ ;
 wire \soc/cpu/_00175_ ;
 wire \soc/cpu/_00176_ ;
 wire \soc/cpu/_00177_ ;
 wire \soc/cpu/_00178_ ;
 wire \soc/cpu/_00179_ ;
 wire \soc/cpu/_00180_ ;
 wire \soc/cpu/_00181_ ;
 wire \soc/cpu/_00182_ ;
 wire \soc/cpu/_00183_ ;
 wire \soc/cpu/_00184_ ;
 wire \soc/cpu/_00185_ ;
 wire \soc/cpu/_00186_ ;
 wire \soc/cpu/_00187_ ;
 wire \soc/cpu/_00188_ ;
 wire \soc/cpu/_00189_ ;
 wire \soc/cpu/_00190_ ;
 wire \soc/cpu/_00191_ ;
 wire \soc/cpu/_00192_ ;
 wire \soc/cpu/_00193_ ;
 wire \soc/cpu/_00194_ ;
 wire \soc/cpu/_00195_ ;
 wire \soc/cpu/_00196_ ;
 wire \soc/cpu/_00197_ ;
 wire \soc/cpu/_00198_ ;
 wire \soc/cpu/_00199_ ;
 wire \soc/cpu/_00200_ ;
 wire \soc/cpu/_00201_ ;
 wire \soc/cpu/_00202_ ;
 wire \soc/cpu/_00203_ ;
 wire \soc/cpu/_00204_ ;
 wire \soc/cpu/_00205_ ;
 wire \soc/cpu/_00206_ ;
 wire \soc/cpu/_00207_ ;
 wire \soc/cpu/_00208_ ;
 wire \soc/cpu/_00209_ ;
 wire \soc/cpu/_00210_ ;
 wire \soc/cpu/_00211_ ;
 wire \soc/cpu/_00212_ ;
 wire \soc/cpu/_00213_ ;
 wire \soc/cpu/_00214_ ;
 wire \soc/cpu/_00215_ ;
 wire \soc/cpu/_00216_ ;
 wire \soc/cpu/_00217_ ;
 wire \soc/cpu/_00218_ ;
 wire \soc/cpu/_00219_ ;
 wire \soc/cpu/_00220_ ;
 wire \soc/cpu/_00221_ ;
 wire \soc/cpu/_00222_ ;
 wire \soc/cpu/_00223_ ;
 wire \soc/cpu/_00224_ ;
 wire \soc/cpu/_00225_ ;
 wire \soc/cpu/_00226_ ;
 wire \soc/cpu/_00227_ ;
 wire \soc/cpu/_00228_ ;
 wire \soc/cpu/_00229_ ;
 wire \soc/cpu/_00230_ ;
 wire \soc/cpu/_00231_ ;
 wire \soc/cpu/_00232_ ;
 wire \soc/cpu/_00233_ ;
 wire \soc/cpu/_00234_ ;
 wire \soc/cpu/_00235_ ;
 wire \soc/cpu/_00236_ ;
 wire \soc/cpu/_00237_ ;
 wire \soc/cpu/_00238_ ;
 wire \soc/cpu/_00239_ ;
 wire \soc/cpu/_00240_ ;
 wire \soc/cpu/_00241_ ;
 wire \soc/cpu/_00242_ ;
 wire \soc/cpu/_00243_ ;
 wire \soc/cpu/_00244_ ;
 wire \soc/cpu/_00245_ ;
 wire \soc/cpu/_00246_ ;
 wire \soc/cpu/_00247_ ;
 wire \soc/cpu/_00248_ ;
 wire \soc/cpu/_00249_ ;
 wire \soc/cpu/_00250_ ;
 wire \soc/cpu/_00251_ ;
 wire \soc/cpu/_00252_ ;
 wire \soc/cpu/_00253_ ;
 wire \soc/cpu/_00254_ ;
 wire \soc/cpu/_00255_ ;
 wire \soc/cpu/_00256_ ;
 wire \soc/cpu/_00257_ ;
 wire \soc/cpu/_00258_ ;
 wire \soc/cpu/_00259_ ;
 wire \soc/cpu/_00260_ ;
 wire \soc/cpu/_00261_ ;
 wire \soc/cpu/_00262_ ;
 wire \soc/cpu/_00263_ ;
 wire \soc/cpu/_00264_ ;
 wire \soc/cpu/_00265_ ;
 wire \soc/cpu/_00266_ ;
 wire \soc/cpu/_00267_ ;
 wire \soc/cpu/_00268_ ;
 wire \soc/cpu/_00269_ ;
 wire \soc/cpu/_00270_ ;
 wire \soc/cpu/_00271_ ;
 wire \soc/cpu/_00272_ ;
 wire \soc/cpu/_00273_ ;
 wire \soc/cpu/_00274_ ;
 wire \soc/cpu/_00275_ ;
 wire \soc/cpu/_00276_ ;
 wire \soc/cpu/_00277_ ;
 wire \soc/cpu/_00278_ ;
 wire \soc/cpu/_00279_ ;
 wire \soc/cpu/_00280_ ;
 wire \soc/cpu/_00281_ ;
 wire \soc/cpu/_00282_ ;
 wire \soc/cpu/_00283_ ;
 wire \soc/cpu/_00284_ ;
 wire \soc/cpu/_00285_ ;
 wire \soc/cpu/_00286_ ;
 wire \soc/cpu/_00287_ ;
 wire \soc/cpu/_00288_ ;
 wire \soc/cpu/_00289_ ;
 wire \soc/cpu/_00290_ ;
 wire \soc/cpu/_00291_ ;
 wire \soc/cpu/_00292_ ;
 wire \soc/cpu/_00293_ ;
 wire \soc/cpu/_00294_ ;
 wire \soc/cpu/_00295_ ;
 wire \soc/cpu/_00296_ ;
 wire \soc/cpu/_00297_ ;
 wire \soc/cpu/_00298_ ;
 wire \soc/cpu/_00299_ ;
 wire \soc/cpu/_00300_ ;
 wire \soc/cpu/_00301_ ;
 wire \soc/cpu/_00302_ ;
 wire \soc/cpu/_00303_ ;
 wire \soc/cpu/_00304_ ;
 wire \soc/cpu/_00305_ ;
 wire \soc/cpu/_00306_ ;
 wire \soc/cpu/_00307_ ;
 wire \soc/cpu/_00308_ ;
 wire \soc/cpu/_00309_ ;
 wire \soc/cpu/_00310_ ;
 wire \soc/cpu/_00311_ ;
 wire \soc/cpu/_00312_ ;
 wire \soc/cpu/_00313_ ;
 wire \soc/cpu/_00314_ ;
 wire \soc/cpu/_00315_ ;
 wire \soc/cpu/_00316_ ;
 wire \soc/cpu/_00317_ ;
 wire \soc/cpu/_00318_ ;
 wire \soc/cpu/_00319_ ;
 wire \soc/cpu/_00320_ ;
 wire \soc/cpu/_00321_ ;
 wire \soc/cpu/_00322_ ;
 wire \soc/cpu/_00323_ ;
 wire \soc/cpu/_00324_ ;
 wire \soc/cpu/_00325_ ;
 wire \soc/cpu/_00326_ ;
 wire \soc/cpu/_00327_ ;
 wire \soc/cpu/_00328_ ;
 wire \soc/cpu/_00329_ ;
 wire \soc/cpu/_00330_ ;
 wire \soc/cpu/_00331_ ;
 wire \soc/cpu/_00332_ ;
 wire \soc/cpu/_00333_ ;
 wire \soc/cpu/_00334_ ;
 wire \soc/cpu/_00335_ ;
 wire \soc/cpu/_00336_ ;
 wire \soc/cpu/_00337_ ;
 wire \soc/cpu/_00338_ ;
 wire \soc/cpu/_00339_ ;
 wire \soc/cpu/_00340_ ;
 wire \soc/cpu/_00341_ ;
 wire \soc/cpu/_00342_ ;
 wire \soc/cpu/_00343_ ;
 wire \soc/cpu/_00344_ ;
 wire \soc/cpu/_00345_ ;
 wire \soc/cpu/_00346_ ;
 wire \soc/cpu/_00347_ ;
 wire \soc/cpu/_00348_ ;
 wire \soc/cpu/_00349_ ;
 wire \soc/cpu/_00350_ ;
 wire \soc/cpu/_00351_ ;
 wire \soc/cpu/_00352_ ;
 wire \soc/cpu/_00353_ ;
 wire \soc/cpu/_00354_ ;
 wire \soc/cpu/_00355_ ;
 wire \soc/cpu/_00356_ ;
 wire \soc/cpu/_00357_ ;
 wire \soc/cpu/_00358_ ;
 wire \soc/cpu/_00359_ ;
 wire \soc/cpu/_00360_ ;
 wire \soc/cpu/_00361_ ;
 wire \soc/cpu/_00362_ ;
 wire \soc/cpu/_00363_ ;
 wire \soc/cpu/_00364_ ;
 wire \soc/cpu/_00365_ ;
 wire \soc/cpu/_00366_ ;
 wire \soc/cpu/_00367_ ;
 wire \soc/cpu/_00368_ ;
 wire \soc/cpu/_00369_ ;
 wire \soc/cpu/_00370_ ;
 wire \soc/cpu/_00371_ ;
 wire \soc/cpu/_00372_ ;
 wire \soc/cpu/_00373_ ;
 wire \soc/cpu/_00374_ ;
 wire \soc/cpu/_00375_ ;
 wire \soc/cpu/_00376_ ;
 wire \soc/cpu/_00377_ ;
 wire \soc/cpu/_00378_ ;
 wire \soc/cpu/_00379_ ;
 wire \soc/cpu/_00380_ ;
 wire \soc/cpu/_00381_ ;
 wire \soc/cpu/_00382_ ;
 wire \soc/cpu/_00383_ ;
 wire \soc/cpu/_00384_ ;
 wire \soc/cpu/_00385_ ;
 wire \soc/cpu/_00386_ ;
 wire \soc/cpu/_00387_ ;
 wire \soc/cpu/_00388_ ;
 wire \soc/cpu/_00389_ ;
 wire \soc/cpu/_00390_ ;
 wire \soc/cpu/_00391_ ;
 wire \soc/cpu/_00392_ ;
 wire \soc/cpu/_00393_ ;
 wire \soc/cpu/_00394_ ;
 wire \soc/cpu/_00395_ ;
 wire \soc/cpu/_00396_ ;
 wire \soc/cpu/_00397_ ;
 wire \soc/cpu/_00398_ ;
 wire \soc/cpu/_00399_ ;
 wire \soc/cpu/_00400_ ;
 wire \soc/cpu/_00401_ ;
 wire \soc/cpu/_00402_ ;
 wire \soc/cpu/_00403_ ;
 wire \soc/cpu/_00404_ ;
 wire \soc/cpu/_00405_ ;
 wire \soc/cpu/_00406_ ;
 wire \soc/cpu/_00407_ ;
 wire \soc/cpu/_00408_ ;
 wire \soc/cpu/_00409_ ;
 wire \soc/cpu/_00410_ ;
 wire \soc/cpu/_00411_ ;
 wire \soc/cpu/_00412_ ;
 wire \soc/cpu/_00413_ ;
 wire \soc/cpu/_00414_ ;
 wire \soc/cpu/_00415_ ;
 wire \soc/cpu/_00416_ ;
 wire \soc/cpu/_00417_ ;
 wire \soc/cpu/_00418_ ;
 wire \soc/cpu/_00419_ ;
 wire \soc/cpu/_00420_ ;
 wire \soc/cpu/_00421_ ;
 wire \soc/cpu/_00422_ ;
 wire \soc/cpu/_00423_ ;
 wire \soc/cpu/_00424_ ;
 wire \soc/cpu/_00425_ ;
 wire \soc/cpu/_00426_ ;
 wire \soc/cpu/_00427_ ;
 wire \soc/cpu/_00428_ ;
 wire \soc/cpu/_00429_ ;
 wire \soc/cpu/_00430_ ;
 wire \soc/cpu/_00431_ ;
 wire \soc/cpu/_00432_ ;
 wire \soc/cpu/_00433_ ;
 wire \soc/cpu/_00434_ ;
 wire \soc/cpu/_00435_ ;
 wire \soc/cpu/_00436_ ;
 wire \soc/cpu/_00437_ ;
 wire \soc/cpu/_00438_ ;
 wire \soc/cpu/_00439_ ;
 wire \soc/cpu/_00440_ ;
 wire \soc/cpu/_00441_ ;
 wire \soc/cpu/_00442_ ;
 wire \soc/cpu/_00443_ ;
 wire \soc/cpu/_00444_ ;
 wire \soc/cpu/_00445_ ;
 wire \soc/cpu/_00446_ ;
 wire \soc/cpu/_00447_ ;
 wire \soc/cpu/_00448_ ;
 wire \soc/cpu/_00449_ ;
 wire \soc/cpu/_00450_ ;
 wire \soc/cpu/_00451_ ;
 wire \soc/cpu/_00452_ ;
 wire \soc/cpu/_00453_ ;
 wire \soc/cpu/_00454_ ;
 wire \soc/cpu/_00455_ ;
 wire \soc/cpu/_00456_ ;
 wire \soc/cpu/_00457_ ;
 wire \soc/cpu/_00458_ ;
 wire \soc/cpu/_00459_ ;
 wire \soc/cpu/_00460_ ;
 wire \soc/cpu/_00461_ ;
 wire \soc/cpu/_00462_ ;
 wire \soc/cpu/_00463_ ;
 wire \soc/cpu/_00464_ ;
 wire \soc/cpu/_00465_ ;
 wire \soc/cpu/_00466_ ;
 wire \soc/cpu/_00467_ ;
 wire \soc/cpu/_00468_ ;
 wire \soc/cpu/_00469_ ;
 wire \soc/cpu/_00470_ ;
 wire \soc/cpu/_00471_ ;
 wire \soc/cpu/_00472_ ;
 wire \soc/cpu/_00473_ ;
 wire \soc/cpu/_00474_ ;
 wire \soc/cpu/_00475_ ;
 wire \soc/cpu/_00476_ ;
 wire \soc/cpu/_00477_ ;
 wire \soc/cpu/_00478_ ;
 wire \soc/cpu/_00479_ ;
 wire \soc/cpu/_00480_ ;
 wire \soc/cpu/_00481_ ;
 wire \soc/cpu/_00482_ ;
 wire \soc/cpu/_00483_ ;
 wire \soc/cpu/_00484_ ;
 wire \soc/cpu/_00485_ ;
 wire \soc/cpu/_00486_ ;
 wire \soc/cpu/_00487_ ;
 wire \soc/cpu/_00488_ ;
 wire \soc/cpu/_00489_ ;
 wire \soc/cpu/_00490_ ;
 wire \soc/cpu/_00491_ ;
 wire \soc/cpu/_00492_ ;
 wire \soc/cpu/_00493_ ;
 wire \soc/cpu/_00494_ ;
 wire \soc/cpu/_00495_ ;
 wire \soc/cpu/_00496_ ;
 wire \soc/cpu/_00497_ ;
 wire \soc/cpu/_00498_ ;
 wire \soc/cpu/_00499_ ;
 wire \soc/cpu/_00500_ ;
 wire \soc/cpu/_00501_ ;
 wire \soc/cpu/_00502_ ;
 wire \soc/cpu/_00503_ ;
 wire \soc/cpu/_00504_ ;
 wire \soc/cpu/_00505_ ;
 wire \soc/cpu/_00506_ ;
 wire \soc/cpu/_00507_ ;
 wire \soc/cpu/_00508_ ;
 wire \soc/cpu/_00509_ ;
 wire \soc/cpu/_00510_ ;
 wire \soc/cpu/_00511_ ;
 wire \soc/cpu/_00512_ ;
 wire \soc/cpu/_00513_ ;
 wire \soc/cpu/_00514_ ;
 wire \soc/cpu/_00515_ ;
 wire \soc/cpu/_00516_ ;
 wire \soc/cpu/_00517_ ;
 wire \soc/cpu/_00518_ ;
 wire \soc/cpu/_00519_ ;
 wire \soc/cpu/_00520_ ;
 wire \soc/cpu/_00521_ ;
 wire \soc/cpu/_00522_ ;
 wire \soc/cpu/_00523_ ;
 wire \soc/cpu/_00524_ ;
 wire \soc/cpu/_00525_ ;
 wire \soc/cpu/_00526_ ;
 wire \soc/cpu/_00527_ ;
 wire \soc/cpu/_00528_ ;
 wire \soc/cpu/_00529_ ;
 wire \soc/cpu/_00530_ ;
 wire \soc/cpu/_00531_ ;
 wire \soc/cpu/_00532_ ;
 wire \soc/cpu/_00533_ ;
 wire \soc/cpu/_00534_ ;
 wire \soc/cpu/_00535_ ;
 wire \soc/cpu/_00536_ ;
 wire \soc/cpu/_00537_ ;
 wire \soc/cpu/_00538_ ;
 wire \soc/cpu/_00539_ ;
 wire \soc/cpu/_00540_ ;
 wire \soc/cpu/_00541_ ;
 wire \soc/cpu/_00542_ ;
 wire \soc/cpu/_00543_ ;
 wire \soc/cpu/_00544_ ;
 wire \soc/cpu/_00545_ ;
 wire \soc/cpu/_00546_ ;
 wire \soc/cpu/_00547_ ;
 wire \soc/cpu/_00548_ ;
 wire \soc/cpu/_00549_ ;
 wire \soc/cpu/_00550_ ;
 wire \soc/cpu/_00551_ ;
 wire \soc/cpu/_00552_ ;
 wire \soc/cpu/_00553_ ;
 wire \soc/cpu/_00554_ ;
 wire \soc/cpu/_00555_ ;
 wire \soc/cpu/_00556_ ;
 wire \soc/cpu/_00557_ ;
 wire \soc/cpu/_00558_ ;
 wire \soc/cpu/_00559_ ;
 wire \soc/cpu/_00560_ ;
 wire \soc/cpu/_00561_ ;
 wire \soc/cpu/_00562_ ;
 wire \soc/cpu/_00563_ ;
 wire \soc/cpu/_00564_ ;
 wire \soc/cpu/_00565_ ;
 wire \soc/cpu/_00566_ ;
 wire \soc/cpu/_00567_ ;
 wire \soc/cpu/_00568_ ;
 wire \soc/cpu/_00569_ ;
 wire \soc/cpu/_00570_ ;
 wire \soc/cpu/_00571_ ;
 wire \soc/cpu/_00572_ ;
 wire \soc/cpu/_00573_ ;
 wire \soc/cpu/_00574_ ;
 wire \soc/cpu/_00575_ ;
 wire \soc/cpu/_00576_ ;
 wire \soc/cpu/_00577_ ;
 wire \soc/cpu/_00578_ ;
 wire \soc/cpu/_00579_ ;
 wire \soc/cpu/_00580_ ;
 wire \soc/cpu/_00581_ ;
 wire \soc/cpu/_00582_ ;
 wire \soc/cpu/_00583_ ;
 wire \soc/cpu/_00584_ ;
 wire \soc/cpu/_00585_ ;
 wire \soc/cpu/_00586_ ;
 wire \soc/cpu/_00587_ ;
 wire \soc/cpu/_00588_ ;
 wire \soc/cpu/_00589_ ;
 wire \soc/cpu/_00590_ ;
 wire \soc/cpu/_00591_ ;
 wire \soc/cpu/_00592_ ;
 wire \soc/cpu/_00593_ ;
 wire \soc/cpu/_00594_ ;
 wire \soc/cpu/_00595_ ;
 wire \soc/cpu/_00596_ ;
 wire \soc/cpu/_00597_ ;
 wire \soc/cpu/_00598_ ;
 wire \soc/cpu/_00599_ ;
 wire \soc/cpu/_00600_ ;
 wire \soc/cpu/_00601_ ;
 wire \soc/cpu/_00602_ ;
 wire \soc/cpu/_00603_ ;
 wire \soc/cpu/_00604_ ;
 wire \soc/cpu/_00605_ ;
 wire \soc/cpu/_00606_ ;
 wire \soc/cpu/_00607_ ;
 wire \soc/cpu/_00608_ ;
 wire \soc/cpu/_00609_ ;
 wire \soc/cpu/_00610_ ;
 wire \soc/cpu/_00611_ ;
 wire \soc/cpu/_00612_ ;
 wire \soc/cpu/_00613_ ;
 wire \soc/cpu/_00614_ ;
 wire \soc/cpu/_00615_ ;
 wire \soc/cpu/_00616_ ;
 wire \soc/cpu/_00617_ ;
 wire \soc/cpu/_00618_ ;
 wire \soc/cpu/_00619_ ;
 wire \soc/cpu/_00620_ ;
 wire \soc/cpu/_00621_ ;
 wire \soc/cpu/_00622_ ;
 wire \soc/cpu/_00623_ ;
 wire \soc/cpu/_00624_ ;
 wire \soc/cpu/_00625_ ;
 wire \soc/cpu/_00626_ ;
 wire \soc/cpu/_00627_ ;
 wire \soc/cpu/_00628_ ;
 wire \soc/cpu/_00629_ ;
 wire \soc/cpu/_00630_ ;
 wire \soc/cpu/_00631_ ;
 wire \soc/cpu/_00632_ ;
 wire \soc/cpu/_00633_ ;
 wire \soc/cpu/_00634_ ;
 wire \soc/cpu/_00635_ ;
 wire \soc/cpu/_00636_ ;
 wire \soc/cpu/_00637_ ;
 wire \soc/cpu/_00638_ ;
 wire \soc/cpu/_00639_ ;
 wire \soc/cpu/_00640_ ;
 wire \soc/cpu/_00641_ ;
 wire \soc/cpu/_00642_ ;
 wire \soc/cpu/_00643_ ;
 wire \soc/cpu/_00644_ ;
 wire \soc/cpu/_00645_ ;
 wire \soc/cpu/_00646_ ;
 wire \soc/cpu/_00647_ ;
 wire \soc/cpu/_00648_ ;
 wire \soc/cpu/_00649_ ;
 wire \soc/cpu/_00650_ ;
 wire \soc/cpu/_00651_ ;
 wire \soc/cpu/_00652_ ;
 wire \soc/cpu/_00653_ ;
 wire \soc/cpu/_00654_ ;
 wire \soc/cpu/_00655_ ;
 wire \soc/cpu/_00656_ ;
 wire \soc/cpu/_00657_ ;
 wire \soc/cpu/_00658_ ;
 wire \soc/cpu/_00659_ ;
 wire \soc/cpu/_00660_ ;
 wire \soc/cpu/_00661_ ;
 wire \soc/cpu/_00662_ ;
 wire \soc/cpu/_00663_ ;
 wire \soc/cpu/_00664_ ;
 wire \soc/cpu/_00665_ ;
 wire \soc/cpu/_00666_ ;
 wire \soc/cpu/_00667_ ;
 wire \soc/cpu/_00668_ ;
 wire \soc/cpu/_00669_ ;
 wire \soc/cpu/_00670_ ;
 wire \soc/cpu/_00671_ ;
 wire \soc/cpu/_00672_ ;
 wire \soc/cpu/_00673_ ;
 wire \soc/cpu/_00674_ ;
 wire \soc/cpu/_00675_ ;
 wire \soc/cpu/_00676_ ;
 wire \soc/cpu/_00677_ ;
 wire \soc/cpu/_00678_ ;
 wire \soc/cpu/_00679_ ;
 wire \soc/cpu/_00680_ ;
 wire \soc/cpu/_00681_ ;
 wire \soc/cpu/_00682_ ;
 wire \soc/cpu/_00683_ ;
 wire \soc/cpu/_00684_ ;
 wire \soc/cpu/_00685_ ;
 wire \soc/cpu/_00686_ ;
 wire \soc/cpu/_00687_ ;
 wire \soc/cpu/_00688_ ;
 wire \soc/cpu/_00689_ ;
 wire \soc/cpu/_00690_ ;
 wire \soc/cpu/_00691_ ;
 wire \soc/cpu/_00692_ ;
 wire \soc/cpu/_00693_ ;
 wire \soc/cpu/_00694_ ;
 wire \soc/cpu/_00695_ ;
 wire \soc/cpu/_00696_ ;
 wire \soc/cpu/_00697_ ;
 wire \soc/cpu/_00698_ ;
 wire \soc/cpu/_00699_ ;
 wire \soc/cpu/_00700_ ;
 wire \soc/cpu/_00701_ ;
 wire \soc/cpu/_00704_ ;
 wire \soc/cpu/_00705_ ;
 wire \soc/cpu/_00707_ ;
 wire \soc/cpu/_00708_ ;
 wire \soc/cpu/_00709_ ;
 wire \soc/cpu/_00711_ ;
 wire \soc/cpu/_00712_ ;
 wire \soc/cpu/_00713_ ;
 wire \soc/cpu/_00714_ ;
 wire \soc/cpu/_00715_ ;
 wire \soc/cpu/_00716_ ;
 wire \soc/cpu/_00718_ ;
 wire \soc/cpu/_00721_ ;
 wire \soc/cpu/_00723_ ;
 wire \soc/cpu/_00724_ ;
 wire \soc/cpu/_00725_ ;
 wire \soc/cpu/_00727_ ;
 wire \soc/cpu/_00728_ ;
 wire \soc/cpu/_00729_ ;
 wire \soc/cpu/_00730_ ;
 wire \soc/cpu/_00732_ ;
 wire \soc/cpu/_00733_ ;
 wire \soc/cpu/_00734_ ;
 wire \soc/cpu/_00735_ ;
 wire \soc/cpu/_00736_ ;
 wire \soc/cpu/_00737_ ;
 wire \soc/cpu/_00738_ ;
 wire \soc/cpu/_00739_ ;
 wire \soc/cpu/_00740_ ;
 wire \soc/cpu/_00741_ ;
 wire \soc/cpu/_00742_ ;
 wire \soc/cpu/_00743_ ;
 wire \soc/cpu/_00744_ ;
 wire \soc/cpu/_00745_ ;
 wire \soc/cpu/_00746_ ;
 wire \soc/cpu/_00747_ ;
 wire \soc/cpu/_00748_ ;
 wire \soc/cpu/_00749_ ;
 wire \soc/cpu/_00750_ ;
 wire \soc/cpu/_00751_ ;
 wire \soc/cpu/_00752_ ;
 wire \soc/cpu/_00753_ ;
 wire \soc/cpu/_00754_ ;
 wire \soc/cpu/_00755_ ;
 wire \soc/cpu/_00756_ ;
 wire \soc/cpu/_00757_ ;
 wire \soc/cpu/_00758_ ;
 wire \soc/cpu/_00759_ ;
 wire \soc/cpu/_00760_ ;
 wire \soc/cpu/_00761_ ;
 wire \soc/cpu/_00762_ ;
 wire \soc/cpu/_00763_ ;
 wire \soc/cpu/_00764_ ;
 wire \soc/cpu/_00765_ ;
 wire \soc/cpu/_00766_ ;
 wire \soc/cpu/_00767_ ;
 wire \soc/cpu/_00768_ ;
 wire \soc/cpu/_00769_ ;
 wire \soc/cpu/_00770_ ;
 wire \soc/cpu/_00771_ ;
 wire \soc/cpu/_00772_ ;
 wire \soc/cpu/_00773_ ;
 wire \soc/cpu/_00774_ ;
 wire \soc/cpu/_00775_ ;
 wire \soc/cpu/_00776_ ;
 wire \soc/cpu/_00777_ ;
 wire \soc/cpu/_00778_ ;
 wire \soc/cpu/_00779_ ;
 wire \soc/cpu/_00780_ ;
 wire \soc/cpu/_00781_ ;
 wire \soc/cpu/_00782_ ;
 wire \soc/cpu/_00783_ ;
 wire \soc/cpu/_00784_ ;
 wire \soc/cpu/_00785_ ;
 wire \soc/cpu/_00786_ ;
 wire \soc/cpu/_00787_ ;
 wire \soc/cpu/_00788_ ;
 wire \soc/cpu/_00789_ ;
 wire \soc/cpu/_00790_ ;
 wire \soc/cpu/_00791_ ;
 wire \soc/cpu/_00795_ ;
 wire \soc/cpu/_00796_ ;
 wire \soc/cpu/_00797_ ;
 wire \soc/cpu/_00800_ ;
 wire \soc/cpu/_00801_ ;
 wire \soc/cpu/_00802_ ;
 wire \soc/cpu/_00803_ ;
 wire \soc/cpu/_00805_ ;
 wire \soc/cpu/_00806_ ;
 wire \soc/cpu/_00807_ ;
 wire \soc/cpu/_00808_ ;
 wire \soc/cpu/_00811_ ;
 wire \soc/cpu/_00812_ ;
 wire \soc/cpu/_00813_ ;
 wire \soc/cpu/_00814_ ;
 wire \soc/cpu/_00815_ ;
 wire \soc/cpu/_00816_ ;
 wire \soc/cpu/_00818_ ;
 wire \soc/cpu/_00822_ ;
 wire \soc/cpu/_00825_ ;
 wire \soc/cpu/_00826_ ;
 wire \soc/cpu/_00827_ ;
 wire \soc/cpu/_00829_ ;
 wire \soc/cpu/_00830_ ;
 wire \soc/cpu/_00831_ ;
 wire \soc/cpu/_00832_ ;
 wire \soc/cpu/_00833_ ;
 wire \soc/cpu/_00834_ ;
 wire \soc/cpu/_00835_ ;
 wire \soc/cpu/_00836_ ;
 wire \soc/cpu/_00837_ ;
 wire \soc/cpu/_00838_ ;
 wire \soc/cpu/_00839_ ;
 wire \soc/cpu/_00840_ ;
 wire \soc/cpu/_00841_ ;
 wire \soc/cpu/_00842_ ;
 wire \soc/cpu/_00843_ ;
 wire \soc/cpu/_00844_ ;
 wire \soc/cpu/_00845_ ;
 wire \soc/cpu/_00846_ ;
 wire \soc/cpu/_00847_ ;
 wire \soc/cpu/_00848_ ;
 wire \soc/cpu/_00849_ ;
 wire \soc/cpu/_00850_ ;
 wire \soc/cpu/_00851_ ;
 wire \soc/cpu/_00852_ ;
 wire \soc/cpu/_00853_ ;
 wire \soc/cpu/_00856_ ;
 wire \soc/cpu/_00857_ ;
 wire \soc/cpu/_00858_ ;
 wire \soc/cpu/_00859_ ;
 wire \soc/cpu/_00861_ ;
 wire \soc/cpu/_00863_ ;
 wire \soc/cpu/_00864_ ;
 wire \soc/cpu/_00865_ ;
 wire \soc/cpu/_00866_ ;
 wire \soc/cpu/_00867_ ;
 wire \soc/cpu/_00868_ ;
 wire \soc/cpu/_00872_ ;
 wire \soc/cpu/_00873_ ;
 wire \soc/cpu/_00874_ ;
 wire \soc/cpu/_00875_ ;
 wire \soc/cpu/_00876_ ;
 wire \soc/cpu/_00877_ ;
 wire \soc/cpu/_00878_ ;
 wire \soc/cpu/_00879_ ;
 wire \soc/cpu/_00880_ ;
 wire \soc/cpu/_00881_ ;
 wire \soc/cpu/_00885_ ;
 wire \soc/cpu/_00886_ ;
 wire \soc/cpu/_00887_ ;
 wire \soc/cpu/_00888_ ;
 wire \soc/cpu/_00889_ ;
 wire \soc/cpu/_00890_ ;
 wire \soc/cpu/_00891_ ;
 wire \soc/cpu/_00892_ ;
 wire \soc/cpu/_00894_ ;
 wire \soc/cpu/_00899_ ;
 wire \soc/cpu/_00900_ ;
 wire \soc/cpu/_00901_ ;
 wire \soc/cpu/_00902_ ;
 wire \soc/cpu/_00903_ ;
 wire \soc/cpu/_00904_ ;
 wire \soc/cpu/_00905_ ;
 wire \soc/cpu/_00906_ ;
 wire \soc/cpu/_00908_ ;
 wire \soc/cpu/_00909_ ;
 wire \soc/cpu/_00910_ ;
 wire \soc/cpu/_00911_ ;
 wire \soc/cpu/_00912_ ;
 wire \soc/cpu/_00914_ ;
 wire \soc/cpu/_00917_ ;
 wire \soc/cpu/_00918_ ;
 wire \soc/cpu/_00919_ ;
 wire \soc/cpu/_00921_ ;
 wire \soc/cpu/_00923_ ;
 wire \soc/cpu/_00924_ ;
 wire \soc/cpu/_00925_ ;
 wire \soc/cpu/_00926_ ;
 wire \soc/cpu/_00928_ ;
 wire \soc/cpu/_00929_ ;
 wire \soc/cpu/_00930_ ;
 wire \soc/cpu/_00931_ ;
 wire \soc/cpu/_00932_ ;
 wire \soc/cpu/_00933_ ;
 wire \soc/cpu/_00934_ ;
 wire \soc/cpu/_00935_ ;
 wire \soc/cpu/_00936_ ;
 wire \soc/cpu/_00937_ ;
 wire \soc/cpu/_00938_ ;
 wire \soc/cpu/_00939_ ;
 wire \soc/cpu/_00940_ ;
 wire \soc/cpu/_00941_ ;
 wire \soc/cpu/_00942_ ;
 wire \soc/cpu/_00943_ ;
 wire \soc/cpu/_00944_ ;
 wire \soc/cpu/_00945_ ;
 wire \soc/cpu/_00946_ ;
 wire \soc/cpu/_00947_ ;
 wire \soc/cpu/_00948_ ;
 wire \soc/cpu/_00950_ ;
 wire \soc/cpu/_00951_ ;
 wire \soc/cpu/_00952_ ;
 wire \soc/cpu/_00953_ ;
 wire \soc/cpu/_00954_ ;
 wire \soc/cpu/_00955_ ;
 wire \soc/cpu/_00956_ ;
 wire \soc/cpu/_00957_ ;
 wire \soc/cpu/_00958_ ;
 wire \soc/cpu/_00960_ ;
 wire \soc/cpu/_00961_ ;
 wire \soc/cpu/_00963_ ;
 wire \soc/cpu/_00964_ ;
 wire \soc/cpu/_00965_ ;
 wire \soc/cpu/_00966_ ;
 wire \soc/cpu/_00969_ ;
 wire \soc/cpu/_00971_ ;
 wire \soc/cpu/_00972_ ;
 wire \soc/cpu/_00973_ ;
 wire \soc/cpu/_00974_ ;
 wire \soc/cpu/_00976_ ;
 wire \soc/cpu/_00979_ ;
 wire \soc/cpu/_00980_ ;
 wire \soc/cpu/_00981_ ;
 wire \soc/cpu/_00982_ ;
 wire \soc/cpu/_00983_ ;
 wire \soc/cpu/_00984_ ;
 wire \soc/cpu/_00985_ ;
 wire \soc/cpu/_00986_ ;
 wire \soc/cpu/_00987_ ;
 wire \soc/cpu/_00989_ ;
 wire \soc/cpu/_00990_ ;
 wire \soc/cpu/_00991_ ;
 wire \soc/cpu/_00992_ ;
 wire \soc/cpu/_00995_ ;
 wire \soc/cpu/_00996_ ;
 wire \soc/cpu/_00997_ ;
 wire \soc/cpu/_00998_ ;
 wire \soc/cpu/_00999_ ;
 wire \soc/cpu/_01000_ ;
 wire \soc/cpu/_01001_ ;
 wire \soc/cpu/_01002_ ;
 wire \soc/cpu/_01003_ ;
 wire \soc/cpu/_01004_ ;
 wire \soc/cpu/_01005_ ;
 wire \soc/cpu/_01006_ ;
 wire \soc/cpu/_01007_ ;
 wire \soc/cpu/_01008_ ;
 wire \soc/cpu/_01009_ ;
 wire \soc/cpu/_01010_ ;
 wire \soc/cpu/_01011_ ;
 wire \soc/cpu/_01012_ ;
 wire \soc/cpu/_01013_ ;
 wire \soc/cpu/_01014_ ;
 wire \soc/cpu/_01015_ ;
 wire \soc/cpu/_01016_ ;
 wire \soc/cpu/_01017_ ;
 wire \soc/cpu/_01018_ ;
 wire \soc/cpu/_01019_ ;
 wire \soc/cpu/_01020_ ;
 wire \soc/cpu/_01021_ ;
 wire \soc/cpu/_01022_ ;
 wire \soc/cpu/_01023_ ;
 wire \soc/cpu/_01024_ ;
 wire \soc/cpu/_01025_ ;
 wire \soc/cpu/_01026_ ;
 wire \soc/cpu/_01027_ ;
 wire \soc/cpu/_01028_ ;
 wire \soc/cpu/_01029_ ;
 wire \soc/cpu/_01030_ ;
 wire \soc/cpu/_01031_ ;
 wire \soc/cpu/_01032_ ;
 wire \soc/cpu/_01033_ ;
 wire \soc/cpu/_01034_ ;
 wire \soc/cpu/_01035_ ;
 wire \soc/cpu/_01036_ ;
 wire \soc/cpu/_01037_ ;
 wire \soc/cpu/_01038_ ;
 wire \soc/cpu/_01039_ ;
 wire \soc/cpu/_01040_ ;
 wire \soc/cpu/_01041_ ;
 wire \soc/cpu/_01042_ ;
 wire \soc/cpu/_01043_ ;
 wire \soc/cpu/_01044_ ;
 wire \soc/cpu/_01045_ ;
 wire \soc/cpu/_01047_ ;
 wire \soc/cpu/_01048_ ;
 wire \soc/cpu/_01050_ ;
 wire \soc/cpu/_01051_ ;
 wire \soc/cpu/_01053_ ;
 wire \soc/cpu/_01054_ ;
 wire \soc/cpu/_01055_ ;
 wire \soc/cpu/_01056_ ;
 wire \soc/cpu/_01057_ ;
 wire \soc/cpu/_01059_ ;
 wire \soc/cpu/_01060_ ;
 wire \soc/cpu/_01061_ ;
 wire \soc/cpu/_01062_ ;
 wire \soc/cpu/_01063_ ;
 wire \soc/cpu/_01064_ ;
 wire \soc/cpu/_01067_ ;
 wire \soc/cpu/_01068_ ;
 wire \soc/cpu/_01069_ ;
 wire \soc/cpu/_01070_ ;
 wire \soc/cpu/_01071_ ;
 wire \soc/cpu/_01072_ ;
 wire \soc/cpu/_01073_ ;
 wire \soc/cpu/_01074_ ;
 wire \soc/cpu/_01075_ ;
 wire \soc/cpu/_01076_ ;
 wire \soc/cpu/_01077_ ;
 wire \soc/cpu/_01078_ ;
 wire \soc/cpu/_01080_ ;
 wire \soc/cpu/_01081_ ;
 wire \soc/cpu/_01082_ ;
 wire \soc/cpu/_01083_ ;
 wire \soc/cpu/_01084_ ;
 wire \soc/cpu/_01085_ ;
 wire \soc/cpu/_01086_ ;
 wire \soc/cpu/_01087_ ;
 wire \soc/cpu/_01088_ ;
 wire \soc/cpu/_01089_ ;
 wire \soc/cpu/_01090_ ;
 wire \soc/cpu/_01091_ ;
 wire \soc/cpu/_01092_ ;
 wire \soc/cpu/_01093_ ;
 wire \soc/cpu/_01094_ ;
 wire \soc/cpu/_01095_ ;
 wire \soc/cpu/_01096_ ;
 wire \soc/cpu/_01097_ ;
 wire \soc/cpu/_01098_ ;
 wire \soc/cpu/_01099_ ;
 wire \soc/cpu/_01100_ ;
 wire \soc/cpu/_01101_ ;
 wire \soc/cpu/_01102_ ;
 wire \soc/cpu/_01103_ ;
 wire \soc/cpu/_01105_ ;
 wire \soc/cpu/_01106_ ;
 wire \soc/cpu/_01107_ ;
 wire \soc/cpu/_01108_ ;
 wire \soc/cpu/_01109_ ;
 wire \soc/cpu/_01110_ ;
 wire \soc/cpu/_01111_ ;
 wire \soc/cpu/_01112_ ;
 wire \soc/cpu/_01113_ ;
 wire \soc/cpu/_01114_ ;
 wire \soc/cpu/_01115_ ;
 wire \soc/cpu/_01116_ ;
 wire \soc/cpu/_01117_ ;
 wire \soc/cpu/_01118_ ;
 wire \soc/cpu/_01120_ ;
 wire \soc/cpu/_01121_ ;
 wire \soc/cpu/_01122_ ;
 wire \soc/cpu/_01123_ ;
 wire \soc/cpu/_01124_ ;
 wire \soc/cpu/_01125_ ;
 wire \soc/cpu/_01126_ ;
 wire \soc/cpu/_01127_ ;
 wire \soc/cpu/_01128_ ;
 wire \soc/cpu/_01129_ ;
 wire \soc/cpu/_01130_ ;
 wire \soc/cpu/_01131_ ;
 wire \soc/cpu/_01132_ ;
 wire \soc/cpu/_01133_ ;
 wire \soc/cpu/_01134_ ;
 wire \soc/cpu/_01135_ ;
 wire \soc/cpu/_01136_ ;
 wire \soc/cpu/_01137_ ;
 wire \soc/cpu/_01138_ ;
 wire \soc/cpu/_01139_ ;
 wire \soc/cpu/_01140_ ;
 wire \soc/cpu/_01141_ ;
 wire \soc/cpu/_01142_ ;
 wire \soc/cpu/_01143_ ;
 wire \soc/cpu/_01144_ ;
 wire \soc/cpu/_01145_ ;
 wire \soc/cpu/_01146_ ;
 wire \soc/cpu/_01147_ ;
 wire \soc/cpu/_01148_ ;
 wire \soc/cpu/_01149_ ;
 wire \soc/cpu/_01150_ ;
 wire \soc/cpu/_01151_ ;
 wire \soc/cpu/_01152_ ;
 wire \soc/cpu/_01153_ ;
 wire \soc/cpu/_01154_ ;
 wire \soc/cpu/_01155_ ;
 wire \soc/cpu/_01156_ ;
 wire \soc/cpu/_01158_ ;
 wire \soc/cpu/_01159_ ;
 wire \soc/cpu/_01160_ ;
 wire \soc/cpu/_01161_ ;
 wire \soc/cpu/_01162_ ;
 wire \soc/cpu/_01163_ ;
 wire \soc/cpu/_01164_ ;
 wire \soc/cpu/_01165_ ;
 wire \soc/cpu/_01166_ ;
 wire \soc/cpu/_01169_ ;
 wire \soc/cpu/_01170_ ;
 wire \soc/cpu/_01171_ ;
 wire \soc/cpu/_01172_ ;
 wire \soc/cpu/_01173_ ;
 wire \soc/cpu/_01174_ ;
 wire \soc/cpu/_01175_ ;
 wire \soc/cpu/_01176_ ;
 wire \soc/cpu/_01177_ ;
 wire \soc/cpu/_01178_ ;
 wire \soc/cpu/_01179_ ;
 wire \soc/cpu/_01180_ ;
 wire \soc/cpu/_01181_ ;
 wire \soc/cpu/_01183_ ;
 wire \soc/cpu/_01185_ ;
 wire \soc/cpu/_01186_ ;
 wire \soc/cpu/_01187_ ;
 wire \soc/cpu/_01188_ ;
 wire \soc/cpu/_01189_ ;
 wire \soc/cpu/_01191_ ;
 wire \soc/cpu/_01192_ ;
 wire \soc/cpu/_01193_ ;
 wire \soc/cpu/_01194_ ;
 wire \soc/cpu/_01195_ ;
 wire \soc/cpu/_01196_ ;
 wire \soc/cpu/_01197_ ;
 wire \soc/cpu/_01198_ ;
 wire \soc/cpu/_01199_ ;
 wire \soc/cpu/_01200_ ;
 wire \soc/cpu/_01201_ ;
 wire \soc/cpu/_01205_ ;
 wire \soc/cpu/_01206_ ;
 wire \soc/cpu/_01207_ ;
 wire \soc/cpu/_01208_ ;
 wire \soc/cpu/_01209_ ;
 wire \soc/cpu/_01210_ ;
 wire \soc/cpu/_01211_ ;
 wire \soc/cpu/_01212_ ;
 wire \soc/cpu/_01213_ ;
 wire \soc/cpu/_01214_ ;
 wire \soc/cpu/_01215_ ;
 wire \soc/cpu/_01217_ ;
 wire \soc/cpu/_01218_ ;
 wire \soc/cpu/_01219_ ;
 wire \soc/cpu/_01220_ ;
 wire \soc/cpu/_01221_ ;
 wire \soc/cpu/_01222_ ;
 wire \soc/cpu/_01223_ ;
 wire \soc/cpu/_01224_ ;
 wire \soc/cpu/_01225_ ;
 wire \soc/cpu/_01226_ ;
 wire \soc/cpu/_01228_ ;
 wire \soc/cpu/_01229_ ;
 wire \soc/cpu/_01230_ ;
 wire \soc/cpu/_01231_ ;
 wire \soc/cpu/_01232_ ;
 wire \soc/cpu/_01233_ ;
 wire \soc/cpu/_01234_ ;
 wire \soc/cpu/_01235_ ;
 wire \soc/cpu/_01236_ ;
 wire \soc/cpu/_01237_ ;
 wire \soc/cpu/_01238_ ;
 wire \soc/cpu/_01239_ ;
 wire \soc/cpu/_01240_ ;
 wire \soc/cpu/_01241_ ;
 wire \soc/cpu/_01242_ ;
 wire \soc/cpu/_01243_ ;
 wire \soc/cpu/_01244_ ;
 wire \soc/cpu/_01245_ ;
 wire \soc/cpu/_01246_ ;
 wire \soc/cpu/_01247_ ;
 wire \soc/cpu/_01248_ ;
 wire \soc/cpu/_01249_ ;
 wire \soc/cpu/_01250_ ;
 wire \soc/cpu/_01251_ ;
 wire \soc/cpu/_01252_ ;
 wire \soc/cpu/_01253_ ;
 wire \soc/cpu/_01254_ ;
 wire \soc/cpu/_01255_ ;
 wire \soc/cpu/_01256_ ;
 wire \soc/cpu/_01257_ ;
 wire \soc/cpu/_01258_ ;
 wire \soc/cpu/_01259_ ;
 wire \soc/cpu/_01260_ ;
 wire \soc/cpu/_01261_ ;
 wire \soc/cpu/_01262_ ;
 wire \soc/cpu/_01263_ ;
 wire \soc/cpu/_01264_ ;
 wire \soc/cpu/_01265_ ;
 wire \soc/cpu/_01266_ ;
 wire \soc/cpu/_01267_ ;
 wire \soc/cpu/_01268_ ;
 wire \soc/cpu/_01270_ ;
 wire \soc/cpu/_01271_ ;
 wire \soc/cpu/_01272_ ;
 wire \soc/cpu/_01273_ ;
 wire \soc/cpu/_01274_ ;
 wire \soc/cpu/_01275_ ;
 wire \soc/cpu/_01276_ ;
 wire \soc/cpu/_01277_ ;
 wire \soc/cpu/_01278_ ;
 wire \soc/cpu/_01279_ ;
 wire \soc/cpu/_01280_ ;
 wire \soc/cpu/_01281_ ;
 wire \soc/cpu/_01282_ ;
 wire \soc/cpu/_01283_ ;
 wire \soc/cpu/_01285_ ;
 wire \soc/cpu/_01286_ ;
 wire \soc/cpu/_01287_ ;
 wire \soc/cpu/_01288_ ;
 wire \soc/cpu/_01289_ ;
 wire \soc/cpu/_01290_ ;
 wire \soc/cpu/_01291_ ;
 wire \soc/cpu/_01293_ ;
 wire \soc/cpu/_01294_ ;
 wire \soc/cpu/_01295_ ;
 wire \soc/cpu/_01296_ ;
 wire \soc/cpu/_01297_ ;
 wire \soc/cpu/_01298_ ;
 wire \soc/cpu/_01300_ ;
 wire \soc/cpu/_01301_ ;
 wire \soc/cpu/_01303_ ;
 wire \soc/cpu/_01304_ ;
 wire \soc/cpu/_01305_ ;
 wire \soc/cpu/_01306_ ;
 wire \soc/cpu/_01308_ ;
 wire \soc/cpu/_01309_ ;
 wire \soc/cpu/_01310_ ;
 wire \soc/cpu/_01311_ ;
 wire \soc/cpu/_01312_ ;
 wire \soc/cpu/_01313_ ;
 wire \soc/cpu/_01314_ ;
 wire \soc/cpu/_01315_ ;
 wire \soc/cpu/_01316_ ;
 wire \soc/cpu/_01317_ ;
 wire \soc/cpu/_01318_ ;
 wire \soc/cpu/_01319_ ;
 wire \soc/cpu/_01320_ ;
 wire \soc/cpu/_01321_ ;
 wire \soc/cpu/_01322_ ;
 wire \soc/cpu/_01323_ ;
 wire \soc/cpu/_01324_ ;
 wire \soc/cpu/_01325_ ;
 wire \soc/cpu/_01326_ ;
 wire \soc/cpu/_01327_ ;
 wire \soc/cpu/_01328_ ;
 wire \soc/cpu/_01329_ ;
 wire \soc/cpu/_01330_ ;
 wire \soc/cpu/_01331_ ;
 wire \soc/cpu/_01333_ ;
 wire \soc/cpu/_01334_ ;
 wire \soc/cpu/_01335_ ;
 wire \soc/cpu/_01336_ ;
 wire \soc/cpu/_01337_ ;
 wire \soc/cpu/_01338_ ;
 wire \soc/cpu/_01339_ ;
 wire \soc/cpu/_01340_ ;
 wire \soc/cpu/_01341_ ;
 wire \soc/cpu/_01342_ ;
 wire \soc/cpu/_01343_ ;
 wire \soc/cpu/_01344_ ;
 wire \soc/cpu/_01345_ ;
 wire \soc/cpu/_01346_ ;
 wire \soc/cpu/_01347_ ;
 wire \soc/cpu/_01348_ ;
 wire \soc/cpu/_01349_ ;
 wire \soc/cpu/_01350_ ;
 wire \soc/cpu/_01351_ ;
 wire \soc/cpu/_01352_ ;
 wire \soc/cpu/_01353_ ;
 wire \soc/cpu/_01354_ ;
 wire \soc/cpu/_01355_ ;
 wire \soc/cpu/_01356_ ;
 wire \soc/cpu/_01357_ ;
 wire \soc/cpu/_01358_ ;
 wire \soc/cpu/_01359_ ;
 wire \soc/cpu/_01360_ ;
 wire \soc/cpu/_01361_ ;
 wire \soc/cpu/_01362_ ;
 wire \soc/cpu/_01363_ ;
 wire \soc/cpu/_01364_ ;
 wire \soc/cpu/_01365_ ;
 wire \soc/cpu/_01366_ ;
 wire \soc/cpu/_01367_ ;
 wire \soc/cpu/_01368_ ;
 wire \soc/cpu/_01369_ ;
 wire \soc/cpu/_01370_ ;
 wire \soc/cpu/_01371_ ;
 wire \soc/cpu/_01372_ ;
 wire \soc/cpu/_01373_ ;
 wire \soc/cpu/_01374_ ;
 wire \soc/cpu/_01375_ ;
 wire \soc/cpu/_01376_ ;
 wire \soc/cpu/_01377_ ;
 wire \soc/cpu/_01378_ ;
 wire \soc/cpu/_01379_ ;
 wire \soc/cpu/_01380_ ;
 wire \soc/cpu/_01381_ ;
 wire \soc/cpu/_01382_ ;
 wire \soc/cpu/_01383_ ;
 wire \soc/cpu/_01384_ ;
 wire \soc/cpu/_01385_ ;
 wire \soc/cpu/_01386_ ;
 wire \soc/cpu/_01387_ ;
 wire \soc/cpu/_01388_ ;
 wire \soc/cpu/_01389_ ;
 wire \soc/cpu/_01390_ ;
 wire \soc/cpu/_01391_ ;
 wire \soc/cpu/_01392_ ;
 wire \soc/cpu/_01393_ ;
 wire \soc/cpu/_01394_ ;
 wire \soc/cpu/_01395_ ;
 wire \soc/cpu/_01396_ ;
 wire \soc/cpu/_01397_ ;
 wire \soc/cpu/_01398_ ;
 wire \soc/cpu/_01399_ ;
 wire \soc/cpu/_01400_ ;
 wire \soc/cpu/_01401_ ;
 wire \soc/cpu/_01402_ ;
 wire \soc/cpu/_01403_ ;
 wire \soc/cpu/_01404_ ;
 wire \soc/cpu/_01405_ ;
 wire \soc/cpu/_01406_ ;
 wire \soc/cpu/_01407_ ;
 wire \soc/cpu/_01408_ ;
 wire \soc/cpu/_01409_ ;
 wire \soc/cpu/_01411_ ;
 wire \soc/cpu/_01412_ ;
 wire \soc/cpu/_01413_ ;
 wire \soc/cpu/_01414_ ;
 wire \soc/cpu/_01415_ ;
 wire \soc/cpu/_01417_ ;
 wire \soc/cpu/_01419_ ;
 wire \soc/cpu/_01420_ ;
 wire \soc/cpu/_01421_ ;
 wire \soc/cpu/_01423_ ;
 wire \soc/cpu/_01424_ ;
 wire \soc/cpu/_01425_ ;
 wire \soc/cpu/_01426_ ;
 wire \soc/cpu/_01427_ ;
 wire \soc/cpu/_01428_ ;
 wire \soc/cpu/_01429_ ;
 wire \soc/cpu/_01431_ ;
 wire \soc/cpu/_01432_ ;
 wire \soc/cpu/_01433_ ;
 wire \soc/cpu/_01435_ ;
 wire \soc/cpu/_01437_ ;
 wire \soc/cpu/_01438_ ;
 wire \soc/cpu/_01439_ ;
 wire \soc/cpu/_01441_ ;
 wire \soc/cpu/_01442_ ;
 wire \soc/cpu/_01443_ ;
 wire \soc/cpu/_01444_ ;
 wire \soc/cpu/_01445_ ;
 wire \soc/cpu/_01448_ ;
 wire \soc/cpu/_01451_ ;
 wire \soc/cpu/_01453_ ;
 wire \soc/cpu/_01454_ ;
 wire \soc/cpu/_01455_ ;
 wire \soc/cpu/_01456_ ;
 wire \soc/cpu/_01458_ ;
 wire \soc/cpu/_01460_ ;
 wire \soc/cpu/_01463_ ;
 wire \soc/cpu/_01464_ ;
 wire \soc/cpu/_01465_ ;
 wire \soc/cpu/_01467_ ;
 wire \soc/cpu/_01470_ ;
 wire \soc/cpu/_01473_ ;
 wire \soc/cpu/_01475_ ;
 wire \soc/cpu/_01476_ ;
 wire \soc/cpu/_01478_ ;
 wire \soc/cpu/_01481_ ;
 wire \soc/cpu/_01482_ ;
 wire \soc/cpu/_01484_ ;
 wire \soc/cpu/_01487_ ;
 wire \soc/cpu/_01488_ ;
 wire \soc/cpu/_01489_ ;
 wire \soc/cpu/_01490_ ;
 wire \soc/cpu/_01492_ ;
 wire \soc/cpu/_01493_ ;
 wire \soc/cpu/_01494_ ;
 wire \soc/cpu/_01496_ ;
 wire \soc/cpu/_01498_ ;
 wire \soc/cpu/_01500_ ;
 wire \soc/cpu/_01501_ ;
 wire \soc/cpu/_01503_ ;
 wire \soc/cpu/_01505_ ;
 wire \soc/cpu/_01506_ ;
 wire \soc/cpu/_01507_ ;
 wire \soc/cpu/_01508_ ;
 wire \soc/cpu/_01510_ ;
 wire \soc/cpu/_01511_ ;
 wire \soc/cpu/_01512_ ;
 wire \soc/cpu/_01513_ ;
 wire \soc/cpu/_01514_ ;
 wire \soc/cpu/_01515_ ;
 wire \soc/cpu/_01516_ ;
 wire \soc/cpu/_01517_ ;
 wire \soc/cpu/_01518_ ;
 wire \soc/cpu/_01519_ ;
 wire \soc/cpu/_01520_ ;
 wire \soc/cpu/_01521_ ;
 wire \soc/cpu/_01522_ ;
 wire \soc/cpu/_01523_ ;
 wire \soc/cpu/_01524_ ;
 wire \soc/cpu/_01525_ ;
 wire \soc/cpu/_01526_ ;
 wire net974;
 wire \soc/cpu/_01528_ ;
 wire \soc/cpu/_01529_ ;
 wire \soc/cpu/_01530_ ;
 wire \soc/cpu/_01531_ ;
 wire \soc/cpu/_01532_ ;
 wire \soc/cpu/_01533_ ;
 wire \soc/cpu/_01534_ ;
 wire \soc/cpu/_01535_ ;
 wire net973;
 wire \soc/cpu/_01537_ ;
 wire \soc/cpu/_01538_ ;
 wire \soc/cpu/_01539_ ;
 wire \soc/cpu/_01540_ ;
 wire \soc/cpu/_01541_ ;
 wire \soc/cpu/_01542_ ;
 wire \soc/cpu/_01543_ ;
 wire \soc/cpu/_01544_ ;
 wire \soc/cpu/_01545_ ;
 wire \soc/cpu/_01546_ ;
 wire \soc/cpu/_01547_ ;
 wire net972;
 wire \soc/cpu/_01549_ ;
 wire net971;
 wire \soc/cpu/_01551_ ;
 wire \soc/cpu/_01552_ ;
 wire net970;
 wire \soc/cpu/_01554_ ;
 wire \soc/cpu/_01555_ ;
 wire \soc/cpu/_01556_ ;
 wire \soc/cpu/_01557_ ;
 wire \soc/cpu/_01558_ ;
 wire \soc/cpu/_01559_ ;
 wire \soc/cpu/_01560_ ;
 wire \soc/cpu/_01561_ ;
 wire \soc/cpu/_01562_ ;
 wire \soc/cpu/_01563_ ;
 wire \soc/cpu/_01564_ ;
 wire \soc/cpu/_01565_ ;
 wire \soc/cpu/_01566_ ;
 wire \soc/cpu/_01567_ ;
 wire \soc/cpu/_01568_ ;
 wire \soc/cpu/_01569_ ;
 wire \soc/cpu/_01570_ ;
 wire \soc/cpu/_01571_ ;
 wire \soc/cpu/_01572_ ;
 wire \soc/cpu/_01573_ ;
 wire \soc/cpu/_01574_ ;
 wire \soc/cpu/_01575_ ;
 wire \soc/cpu/_01576_ ;
 wire \soc/cpu/_01577_ ;
 wire \soc/cpu/_01578_ ;
 wire \soc/cpu/_01579_ ;
 wire \soc/cpu/_01580_ ;
 wire \soc/cpu/_01581_ ;
 wire \soc/cpu/_01582_ ;
 wire \soc/cpu/_01583_ ;
 wire \soc/cpu/_01584_ ;
 wire \soc/cpu/_01585_ ;
 wire \soc/cpu/_01586_ ;
 wire \soc/cpu/_01587_ ;
 wire \soc/cpu/_01588_ ;
 wire net969;
 wire \soc/cpu/_01590_ ;
 wire \soc/cpu/_01591_ ;
 wire \soc/cpu/_01592_ ;
 wire \soc/cpu/_01593_ ;
 wire \soc/cpu/_01594_ ;
 wire \soc/cpu/_01595_ ;
 wire \soc/cpu/_01596_ ;
 wire \soc/cpu/_01597_ ;
 wire \soc/cpu/_01598_ ;
 wire \soc/cpu/_01599_ ;
 wire net968;
 wire \soc/cpu/_01601_ ;
 wire \soc/cpu/_01602_ ;
 wire net967;
 wire \soc/cpu/_01604_ ;
 wire net966;
 wire \soc/cpu/_01606_ ;
 wire \soc/cpu/_01607_ ;
 wire \soc/cpu/_01608_ ;
 wire \soc/cpu/_01609_ ;
 wire \soc/cpu/_01610_ ;
 wire \soc/cpu/_01611_ ;
 wire \soc/cpu/_01612_ ;
 wire net965;
 wire \soc/cpu/_01614_ ;
 wire net964;
 wire \soc/cpu/_01616_ ;
 wire net963;
 wire \soc/cpu/_01618_ ;
 wire \soc/cpu/_01619_ ;
 wire \soc/cpu/_01620_ ;
 wire net962;
 wire \soc/cpu/_01622_ ;
 wire \soc/cpu/_01623_ ;
 wire \soc/cpu/_01624_ ;
 wire \soc/cpu/_01625_ ;
 wire \soc/cpu/_01626_ ;
 wire net961;
 wire \soc/cpu/_01628_ ;
 wire \soc/cpu/_01629_ ;
 wire \soc/cpu/_01630_ ;
 wire \soc/cpu/_01631_ ;
 wire net960;
 wire \soc/cpu/_01633_ ;
 wire \soc/cpu/_01634_ ;
 wire \soc/cpu/_01635_ ;
 wire \soc/cpu/_01636_ ;
 wire \soc/cpu/_01637_ ;
 wire \soc/cpu/_01638_ ;
 wire \soc/cpu/_01639_ ;
 wire \soc/cpu/_01640_ ;
 wire \soc/cpu/_01641_ ;
 wire net959;
 wire \soc/cpu/_01643_ ;
 wire \soc/cpu/_01644_ ;
 wire \soc/cpu/_01645_ ;
 wire \soc/cpu/_01646_ ;
 wire \soc/cpu/_01647_ ;
 wire \soc/cpu/_01648_ ;
 wire \soc/cpu/_01649_ ;
 wire net958;
 wire \soc/cpu/_01651_ ;
 wire net957;
 wire \soc/cpu/_01653_ ;
 wire \soc/cpu/_01654_ ;
 wire \soc/cpu/_01655_ ;
 wire \soc/cpu/_01656_ ;
 wire \soc/cpu/_01657_ ;
 wire net956;
 wire \soc/cpu/_01659_ ;
 wire \soc/cpu/_01660_ ;
 wire \soc/cpu/_01661_ ;
 wire \soc/cpu/_01662_ ;
 wire \soc/cpu/_01663_ ;
 wire \soc/cpu/_01664_ ;
 wire \soc/cpu/_01665_ ;
 wire \soc/cpu/_01666_ ;
 wire \soc/cpu/_01667_ ;
 wire \soc/cpu/_01668_ ;
 wire \soc/cpu/_01669_ ;
 wire \soc/cpu/_01670_ ;
 wire \soc/cpu/_01671_ ;
 wire \soc/cpu/_01672_ ;
 wire \soc/cpu/_01673_ ;
 wire \soc/cpu/_01674_ ;
 wire \soc/cpu/_01675_ ;
 wire \soc/cpu/_01676_ ;
 wire \soc/cpu/_01677_ ;
 wire net955;
 wire \soc/cpu/_01679_ ;
 wire \soc/cpu/_01680_ ;
 wire \soc/cpu/_01681_ ;
 wire net954;
 wire \soc/cpu/_01683_ ;
 wire \soc/cpu/_01684_ ;
 wire \soc/cpu/_01685_ ;
 wire \soc/cpu/_01686_ ;
 wire \soc/cpu/_01687_ ;
 wire \soc/cpu/_01688_ ;
 wire \soc/cpu/_01689_ ;
 wire \soc/cpu/_01690_ ;
 wire \soc/cpu/_01691_ ;
 wire net953;
 wire \soc/cpu/_01693_ ;
 wire \soc/cpu/_01694_ ;
 wire \soc/cpu/_01695_ ;
 wire \soc/cpu/_01696_ ;
 wire \soc/cpu/_01697_ ;
 wire net952;
 wire \soc/cpu/_01699_ ;
 wire \soc/cpu/_01700_ ;
 wire \soc/cpu/_01701_ ;
 wire \soc/cpu/_01702_ ;
 wire \soc/cpu/_01703_ ;
 wire \soc/cpu/_01704_ ;
 wire \soc/cpu/_01705_ ;
 wire \soc/cpu/_01706_ ;
 wire net951;
 wire \soc/cpu/_01708_ ;
 wire \soc/cpu/_01709_ ;
 wire \soc/cpu/_01710_ ;
 wire net950;
 wire \soc/cpu/_01712_ ;
 wire \soc/cpu/_01713_ ;
 wire \soc/cpu/_01714_ ;
 wire \soc/cpu/_01715_ ;
 wire net949;
 wire \soc/cpu/_01717_ ;
 wire \soc/cpu/_01718_ ;
 wire \soc/cpu/_01719_ ;
 wire \soc/cpu/_01720_ ;
 wire \soc/cpu/_01721_ ;
 wire \soc/cpu/_01722_ ;
 wire net948;
 wire \soc/cpu/_01724_ ;
 wire \soc/cpu/_01725_ ;
 wire \soc/cpu/_01726_ ;
 wire net947;
 wire \soc/cpu/_01728_ ;
 wire \soc/cpu/_01729_ ;
 wire net946;
 wire \soc/cpu/_01731_ ;
 wire \soc/cpu/_01732_ ;
 wire \soc/cpu/_01733_ ;
 wire net945;
 wire \soc/cpu/_01735_ ;
 wire \soc/cpu/_01736_ ;
 wire \soc/cpu/_01737_ ;
 wire \soc/cpu/_01738_ ;
 wire \soc/cpu/_01739_ ;
 wire \soc/cpu/_01740_ ;
 wire net944;
 wire \soc/cpu/_01742_ ;
 wire \soc/cpu/_01743_ ;
 wire \soc/cpu/_01744_ ;
 wire net943;
 wire \soc/cpu/_01746_ ;
 wire \soc/cpu/_01747_ ;
 wire \soc/cpu/_01748_ ;
 wire \soc/cpu/_01749_ ;
 wire \soc/cpu/_01750_ ;
 wire \soc/cpu/_01751_ ;
 wire \soc/cpu/_01752_ ;
 wire net942;
 wire net941;
 wire \soc/cpu/_01755_ ;
 wire \soc/cpu/_01756_ ;
 wire net940;
 wire net939;
 wire \soc/cpu/_01759_ ;
 wire \soc/cpu/_01760_ ;
 wire net938;
 wire \soc/cpu/_01762_ ;
 wire \soc/cpu/_01763_ ;
 wire \soc/cpu/_01764_ ;
 wire net937;
 wire net936;
 wire \soc/cpu/_01767_ ;
 wire \soc/cpu/_01768_ ;
 wire \soc/cpu/_01769_ ;
 wire \soc/cpu/_01770_ ;
 wire \soc/cpu/_01771_ ;
 wire \soc/cpu/_01772_ ;
 wire \soc/cpu/_01773_ ;
 wire \soc/cpu/_01774_ ;
 wire \soc/cpu/_01775_ ;
 wire \soc/cpu/_01776_ ;
 wire \soc/cpu/_01777_ ;
 wire \soc/cpu/_01778_ ;
 wire \soc/cpu/_01779_ ;
 wire net935;
 wire \soc/cpu/_01781_ ;
 wire \soc/cpu/_01782_ ;
 wire \soc/cpu/_01783_ ;
 wire \soc/cpu/_01784_ ;
 wire \soc/cpu/_01785_ ;
 wire \soc/cpu/_01786_ ;
 wire \soc/cpu/_01787_ ;
 wire \soc/cpu/_01788_ ;
 wire \soc/cpu/_01789_ ;
 wire \soc/cpu/_01790_ ;
 wire net934;
 wire \soc/cpu/_01792_ ;
 wire net933;
 wire \soc/cpu/_01794_ ;
 wire \soc/cpu/_01795_ ;
 wire \soc/cpu/_01796_ ;
 wire \soc/cpu/_01797_ ;
 wire net932;
 wire \soc/cpu/_01799_ ;
 wire \soc/cpu/_01800_ ;
 wire net931;
 wire \soc/cpu/_01802_ ;
 wire net930;
 wire \soc/cpu/_01804_ ;
 wire \soc/cpu/_01805_ ;
 wire \soc/cpu/_01806_ ;
 wire \soc/cpu/_01807_ ;
 wire \soc/cpu/_01808_ ;
 wire \soc/cpu/_01809_ ;
 wire \soc/cpu/_01810_ ;
 wire \soc/cpu/_01811_ ;
 wire \soc/cpu/_01812_ ;
 wire \soc/cpu/_01813_ ;
 wire \soc/cpu/_01814_ ;
 wire \soc/cpu/_01815_ ;
 wire \soc/cpu/_01816_ ;
 wire \soc/cpu/_01817_ ;
 wire \soc/cpu/_01818_ ;
 wire \soc/cpu/_01819_ ;
 wire \soc/cpu/_01820_ ;
 wire \soc/cpu/_01821_ ;
 wire \soc/cpu/_01822_ ;
 wire \soc/cpu/_01823_ ;
 wire \soc/cpu/_01824_ ;
 wire \soc/cpu/_01825_ ;
 wire \soc/cpu/_01826_ ;
 wire \soc/cpu/_01827_ ;
 wire \soc/cpu/_01828_ ;
 wire \soc/cpu/_01829_ ;
 wire net929;
 wire \soc/cpu/_01831_ ;
 wire \soc/cpu/_01832_ ;
 wire \soc/cpu/_01833_ ;
 wire \soc/cpu/_01834_ ;
 wire \soc/cpu/_01835_ ;
 wire \soc/cpu/_01836_ ;
 wire \soc/cpu/_01837_ ;
 wire \soc/cpu/_01838_ ;
 wire \soc/cpu/_01839_ ;
 wire \soc/cpu/_01840_ ;
 wire \soc/cpu/_01841_ ;
 wire \soc/cpu/_01842_ ;
 wire \soc/cpu/_01843_ ;
 wire \soc/cpu/_01844_ ;
 wire \soc/cpu/_01845_ ;
 wire \soc/cpu/_01846_ ;
 wire \soc/cpu/_01847_ ;
 wire \soc/cpu/_01848_ ;
 wire \soc/cpu/_01849_ ;
 wire \soc/cpu/_01850_ ;
 wire \soc/cpu/_01851_ ;
 wire \soc/cpu/_01852_ ;
 wire \soc/cpu/_01853_ ;
 wire \soc/cpu/_01854_ ;
 wire \soc/cpu/_01855_ ;
 wire \soc/cpu/_01856_ ;
 wire \soc/cpu/_01857_ ;
 wire \soc/cpu/_01858_ ;
 wire \soc/cpu/_01859_ ;
 wire \soc/cpu/_01860_ ;
 wire \soc/cpu/_01861_ ;
 wire \soc/cpu/_01862_ ;
 wire \soc/cpu/_01863_ ;
 wire \soc/cpu/_01864_ ;
 wire \soc/cpu/_01865_ ;
 wire \soc/cpu/_01866_ ;
 wire \soc/cpu/_01867_ ;
 wire \soc/cpu/_01868_ ;
 wire \soc/cpu/_01869_ ;
 wire \soc/cpu/_01870_ ;
 wire \soc/cpu/_01871_ ;
 wire \soc/cpu/_01872_ ;
 wire \soc/cpu/_01873_ ;
 wire \soc/cpu/_01874_ ;
 wire \soc/cpu/_01875_ ;
 wire \soc/cpu/_01876_ ;
 wire \soc/cpu/_01877_ ;
 wire \soc/cpu/_01878_ ;
 wire \soc/cpu/_01879_ ;
 wire \soc/cpu/_01880_ ;
 wire \soc/cpu/_01881_ ;
 wire \soc/cpu/_01882_ ;
 wire \soc/cpu/_01883_ ;
 wire \soc/cpu/_01884_ ;
 wire \soc/cpu/_01885_ ;
 wire \soc/cpu/_01886_ ;
 wire \soc/cpu/_01887_ ;
 wire \soc/cpu/_01888_ ;
 wire \soc/cpu/_01889_ ;
 wire \soc/cpu/_01890_ ;
 wire \soc/cpu/_01891_ ;
 wire \soc/cpu/_01892_ ;
 wire \soc/cpu/_01893_ ;
 wire \soc/cpu/_01894_ ;
 wire \soc/cpu/_01895_ ;
 wire \soc/cpu/_01896_ ;
 wire \soc/cpu/_01897_ ;
 wire \soc/cpu/_01898_ ;
 wire \soc/cpu/_01899_ ;
 wire \soc/cpu/_01900_ ;
 wire \soc/cpu/_01901_ ;
 wire \soc/cpu/_01902_ ;
 wire \soc/cpu/_01903_ ;
 wire \soc/cpu/_01904_ ;
 wire \soc/cpu/_01905_ ;
 wire \soc/cpu/_01906_ ;
 wire \soc/cpu/_01907_ ;
 wire \soc/cpu/_01908_ ;
 wire \soc/cpu/_01909_ ;
 wire \soc/cpu/_01910_ ;
 wire \soc/cpu/_01911_ ;
 wire \soc/cpu/_01912_ ;
 wire \soc/cpu/_01913_ ;
 wire \soc/cpu/_01914_ ;
 wire \soc/cpu/_01915_ ;
 wire \soc/cpu/_01916_ ;
 wire \soc/cpu/_01917_ ;
 wire \soc/cpu/_01918_ ;
 wire \soc/cpu/_01919_ ;
 wire \soc/cpu/_01920_ ;
 wire \soc/cpu/_01921_ ;
 wire \soc/cpu/_01922_ ;
 wire \soc/cpu/_01923_ ;
 wire \soc/cpu/_01924_ ;
 wire \soc/cpu/_01925_ ;
 wire \soc/cpu/_01926_ ;
 wire \soc/cpu/_01927_ ;
 wire \soc/cpu/_01928_ ;
 wire \soc/cpu/_01929_ ;
 wire \soc/cpu/_01930_ ;
 wire \soc/cpu/_01931_ ;
 wire \soc/cpu/_01932_ ;
 wire \soc/cpu/_01933_ ;
 wire \soc/cpu/_01934_ ;
 wire \soc/cpu/_01935_ ;
 wire \soc/cpu/_01936_ ;
 wire \soc/cpu/_01937_ ;
 wire \soc/cpu/_01938_ ;
 wire \soc/cpu/_01939_ ;
 wire \soc/cpu/_01940_ ;
 wire \soc/cpu/_01941_ ;
 wire \soc/cpu/_01942_ ;
 wire \soc/cpu/_01943_ ;
 wire \soc/cpu/_01944_ ;
 wire \soc/cpu/_01945_ ;
 wire \soc/cpu/_01946_ ;
 wire \soc/cpu/_01947_ ;
 wire \soc/cpu/_01948_ ;
 wire \soc/cpu/_01949_ ;
 wire \soc/cpu/_01950_ ;
 wire \soc/cpu/_01951_ ;
 wire \soc/cpu/_01952_ ;
 wire \soc/cpu/_01953_ ;
 wire \soc/cpu/_01954_ ;
 wire \soc/cpu/_01955_ ;
 wire \soc/cpu/_01956_ ;
 wire \soc/cpu/_01957_ ;
 wire \soc/cpu/_01958_ ;
 wire \soc/cpu/_01959_ ;
 wire \soc/cpu/_01960_ ;
 wire \soc/cpu/_01961_ ;
 wire \soc/cpu/_01962_ ;
 wire \soc/cpu/_01963_ ;
 wire \soc/cpu/_01964_ ;
 wire \soc/cpu/_01965_ ;
 wire \soc/cpu/_01966_ ;
 wire \soc/cpu/_01967_ ;
 wire \soc/cpu/_01968_ ;
 wire \soc/cpu/_01969_ ;
 wire \soc/cpu/_01970_ ;
 wire \soc/cpu/_01971_ ;
 wire \soc/cpu/_01972_ ;
 wire \soc/cpu/_01973_ ;
 wire \soc/cpu/_01974_ ;
 wire \soc/cpu/_01975_ ;
 wire \soc/cpu/_01976_ ;
 wire \soc/cpu/_01977_ ;
 wire \soc/cpu/_01978_ ;
 wire \soc/cpu/_01979_ ;
 wire \soc/cpu/_01980_ ;
 wire \soc/cpu/_01981_ ;
 wire \soc/cpu/_01982_ ;
 wire \soc/cpu/_01983_ ;
 wire \soc/cpu/_01984_ ;
 wire \soc/cpu/_01985_ ;
 wire \soc/cpu/_01986_ ;
 wire \soc/cpu/_01987_ ;
 wire \soc/cpu/_01988_ ;
 wire \soc/cpu/_01989_ ;
 wire \soc/cpu/_01990_ ;
 wire \soc/cpu/_01991_ ;
 wire \soc/cpu/_01992_ ;
 wire \soc/cpu/_01993_ ;
 wire \soc/cpu/_01994_ ;
 wire \soc/cpu/_01995_ ;
 wire \soc/cpu/_01996_ ;
 wire \soc/cpu/_01997_ ;
 wire \soc/cpu/_01998_ ;
 wire \soc/cpu/_01999_ ;
 wire \soc/cpu/_02000_ ;
 wire \soc/cpu/_02001_ ;
 wire \soc/cpu/_02002_ ;
 wire \soc/cpu/_02003_ ;
 wire \soc/cpu/_02004_ ;
 wire \soc/cpu/_02005_ ;
 wire \soc/cpu/_02006_ ;
 wire \soc/cpu/_02007_ ;
 wire \soc/cpu/_02008_ ;
 wire \soc/cpu/_02009_ ;
 wire \soc/cpu/_02010_ ;
 wire \soc/cpu/_02011_ ;
 wire \soc/cpu/_02012_ ;
 wire \soc/cpu/_02013_ ;
 wire \soc/cpu/_02014_ ;
 wire \soc/cpu/_02015_ ;
 wire \soc/cpu/_02016_ ;
 wire \soc/cpu/_02017_ ;
 wire \soc/cpu/_02018_ ;
 wire \soc/cpu/_02019_ ;
 wire \soc/cpu/_02020_ ;
 wire \soc/cpu/_02021_ ;
 wire \soc/cpu/_02022_ ;
 wire \soc/cpu/_02023_ ;
 wire \soc/cpu/_02024_ ;
 wire \soc/cpu/_02025_ ;
 wire \soc/cpu/_02026_ ;
 wire \soc/cpu/_02027_ ;
 wire \soc/cpu/_02028_ ;
 wire \soc/cpu/_02029_ ;
 wire \soc/cpu/_02030_ ;
 wire \soc/cpu/_02031_ ;
 wire \soc/cpu/_02032_ ;
 wire \soc/cpu/_02033_ ;
 wire \soc/cpu/_02034_ ;
 wire \soc/cpu/_02035_ ;
 wire \soc/cpu/_02036_ ;
 wire \soc/cpu/_02037_ ;
 wire \soc/cpu/_02038_ ;
 wire \soc/cpu/_02039_ ;
 wire \soc/cpu/_02040_ ;
 wire \soc/cpu/_02041_ ;
 wire \soc/cpu/_02042_ ;
 wire \soc/cpu/_02043_ ;
 wire \soc/cpu/_02044_ ;
 wire \soc/cpu/_02045_ ;
 wire \soc/cpu/_02046_ ;
 wire \soc/cpu/_02047_ ;
 wire \soc/cpu/_02048_ ;
 wire \soc/cpu/_02049_ ;
 wire \soc/cpu/_02050_ ;
 wire \soc/cpu/_02051_ ;
 wire \soc/cpu/_02052_ ;
 wire \soc/cpu/_02053_ ;
 wire \soc/cpu/_02054_ ;
 wire \soc/cpu/_02055_ ;
 wire \soc/cpu/_02056_ ;
 wire \soc/cpu/_02057_ ;
 wire \soc/cpu/_02058_ ;
 wire \soc/cpu/_02059_ ;
 wire \soc/cpu/_02060_ ;
 wire \soc/cpu/_02061_ ;
 wire \soc/cpu/_02062_ ;
 wire \soc/cpu/_02063_ ;
 wire \soc/cpu/_02064_ ;
 wire \soc/cpu/_02065_ ;
 wire \soc/cpu/_02066_ ;
 wire \soc/cpu/_02067_ ;
 wire \soc/cpu/_02068_ ;
 wire \soc/cpu/_02069_ ;
 wire \soc/cpu/_02070_ ;
 wire \soc/cpu/_02071_ ;
 wire \soc/cpu/_02072_ ;
 wire \soc/cpu/_02073_ ;
 wire \soc/cpu/_02074_ ;
 wire \soc/cpu/_02075_ ;
 wire \soc/cpu/_02076_ ;
 wire \soc/cpu/_02077_ ;
 wire \soc/cpu/_02078_ ;
 wire \soc/cpu/_02079_ ;
 wire \soc/cpu/_02080_ ;
 wire \soc/cpu/_02081_ ;
 wire \soc/cpu/_02082_ ;
 wire \soc/cpu/_02083_ ;
 wire \soc/cpu/_02084_ ;
 wire \soc/cpu/_02085_ ;
 wire \soc/cpu/_02086_ ;
 wire \soc/cpu/_02087_ ;
 wire \soc/cpu/_02088_ ;
 wire \soc/cpu/_02089_ ;
 wire \soc/cpu/_02090_ ;
 wire \soc/cpu/_02091_ ;
 wire \soc/cpu/_02092_ ;
 wire \soc/cpu/_02093_ ;
 wire \soc/cpu/_02094_ ;
 wire \soc/cpu/_02095_ ;
 wire \soc/cpu/_02096_ ;
 wire \soc/cpu/_02097_ ;
 wire \soc/cpu/_02098_ ;
 wire \soc/cpu/_02099_ ;
 wire \soc/cpu/_02100_ ;
 wire \soc/cpu/_02101_ ;
 wire \soc/cpu/_02102_ ;
 wire net928;
 wire net927;
 wire net926;
 wire net925;
 wire \soc/cpu/_02107_ ;
 wire \soc/cpu/_02108_ ;
 wire \soc/cpu/_02109_ ;
 wire net924;
 wire \soc/cpu/_02111_ ;
 wire \soc/cpu/_02112_ ;
 wire net923;
 wire net922;
 wire \soc/cpu/_02115_ ;
 wire net921;
 wire \soc/cpu/_02117_ ;
 wire \soc/cpu/_02118_ ;
 wire \soc/cpu/_02119_ ;
 wire \soc/cpu/_02120_ ;
 wire net920;
 wire net919;
 wire \soc/cpu/_02123_ ;
 wire \soc/cpu/_02124_ ;
 wire \soc/cpu/_02125_ ;
 wire net918;
 wire \soc/cpu/_02127_ ;
 wire net917;
 wire \soc/cpu/_02129_ ;
 wire \soc/cpu/_02130_ ;
 wire net916;
 wire \soc/cpu/_02132_ ;
 wire \soc/cpu/_02133_ ;
 wire \soc/cpu/_02134_ ;
 wire \soc/cpu/_02135_ ;
 wire \soc/cpu/_02136_ ;
 wire \soc/cpu/_02137_ ;
 wire \soc/cpu/_02138_ ;
 wire \soc/cpu/_02139_ ;
 wire \soc/cpu/_02140_ ;
 wire \soc/cpu/_02141_ ;
 wire \soc/cpu/_02142_ ;
 wire \soc/cpu/_02143_ ;
 wire \soc/cpu/_02144_ ;
 wire \soc/cpu/_02145_ ;
 wire \soc/cpu/_02146_ ;
 wire \soc/cpu/_02147_ ;
 wire \soc/cpu/_02148_ ;
 wire net915;
 wire net914;
 wire net913;
 wire \soc/cpu/_02152_ ;
 wire \soc/cpu/_02153_ ;
 wire \soc/cpu/_02154_ ;
 wire net912;
 wire \soc/cpu/_02156_ ;
 wire \soc/cpu/_02157_ ;
 wire \soc/cpu/_02158_ ;
 wire \soc/cpu/_02159_ ;
 wire \soc/cpu/_02160_ ;
 wire \soc/cpu/_02161_ ;
 wire \soc/cpu/_02162_ ;
 wire \soc/cpu/_02163_ ;
 wire \soc/cpu/_02164_ ;
 wire \soc/cpu/_02165_ ;
 wire \soc/cpu/_02166_ ;
 wire \soc/cpu/_02167_ ;
 wire \soc/cpu/_02168_ ;
 wire net911;
 wire \soc/cpu/_02170_ ;
 wire \soc/cpu/_02171_ ;
 wire \soc/cpu/_02172_ ;
 wire \soc/cpu/_02173_ ;
 wire \soc/cpu/_02174_ ;
 wire \soc/cpu/_02175_ ;
 wire \soc/cpu/_02176_ ;
 wire \soc/cpu/_02177_ ;
 wire \soc/cpu/_02178_ ;
 wire \soc/cpu/_02179_ ;
 wire \soc/cpu/_02180_ ;
 wire \soc/cpu/_02181_ ;
 wire \soc/cpu/_02182_ ;
 wire \soc/cpu/_02183_ ;
 wire \soc/cpu/_02184_ ;
 wire \soc/cpu/_02185_ ;
 wire \soc/cpu/_02186_ ;
 wire \soc/cpu/_02187_ ;
 wire \soc/cpu/_02188_ ;
 wire \soc/cpu/_02189_ ;
 wire \soc/cpu/_02190_ ;
 wire \soc/cpu/_02191_ ;
 wire \soc/cpu/_02192_ ;
 wire \soc/cpu/_02193_ ;
 wire \soc/cpu/_02194_ ;
 wire \soc/cpu/_02195_ ;
 wire \soc/cpu/_02196_ ;
 wire \soc/cpu/_02197_ ;
 wire \soc/cpu/_02198_ ;
 wire \soc/cpu/_02199_ ;
 wire \soc/cpu/_02200_ ;
 wire \soc/cpu/_02201_ ;
 wire \soc/cpu/_02202_ ;
 wire \soc/cpu/_02203_ ;
 wire \soc/cpu/_02204_ ;
 wire \soc/cpu/_02205_ ;
 wire \soc/cpu/_02206_ ;
 wire \soc/cpu/_02207_ ;
 wire \soc/cpu/_02208_ ;
 wire \soc/cpu/_02209_ ;
 wire \soc/cpu/_02210_ ;
 wire \soc/cpu/_02211_ ;
 wire \soc/cpu/_02212_ ;
 wire \soc/cpu/_02213_ ;
 wire \soc/cpu/_02214_ ;
 wire \soc/cpu/_02215_ ;
 wire \soc/cpu/_02216_ ;
 wire \soc/cpu/_02217_ ;
 wire \soc/cpu/_02218_ ;
 wire \soc/cpu/_02219_ ;
 wire \soc/cpu/_02220_ ;
 wire \soc/cpu/_02221_ ;
 wire \soc/cpu/_02222_ ;
 wire \soc/cpu/_02223_ ;
 wire \soc/cpu/_02224_ ;
 wire \soc/cpu/_02225_ ;
 wire \soc/cpu/_02226_ ;
 wire \soc/cpu/_02227_ ;
 wire \soc/cpu/_02228_ ;
 wire \soc/cpu/_02229_ ;
 wire \soc/cpu/_02230_ ;
 wire \soc/cpu/_02231_ ;
 wire \soc/cpu/_02232_ ;
 wire \soc/cpu/_02233_ ;
 wire \soc/cpu/_02234_ ;
 wire \soc/cpu/_02235_ ;
 wire \soc/cpu/_02236_ ;
 wire \soc/cpu/_02237_ ;
 wire \soc/cpu/_02238_ ;
 wire \soc/cpu/_02239_ ;
 wire \soc/cpu/_02240_ ;
 wire \soc/cpu/_02241_ ;
 wire \soc/cpu/_02242_ ;
 wire \soc/cpu/_02243_ ;
 wire \soc/cpu/_02244_ ;
 wire \soc/cpu/_02245_ ;
 wire \soc/cpu/_02246_ ;
 wire \soc/cpu/_02247_ ;
 wire \soc/cpu/_02248_ ;
 wire \soc/cpu/_02249_ ;
 wire \soc/cpu/_02250_ ;
 wire \soc/cpu/_02251_ ;
 wire \soc/cpu/_02252_ ;
 wire \soc/cpu/_02253_ ;
 wire \soc/cpu/_02254_ ;
 wire \soc/cpu/_02255_ ;
 wire \soc/cpu/_02256_ ;
 wire \soc/cpu/_02257_ ;
 wire \soc/cpu/_02258_ ;
 wire \soc/cpu/_02259_ ;
 wire \soc/cpu/_02260_ ;
 wire \soc/cpu/_02261_ ;
 wire \soc/cpu/_02262_ ;
 wire \soc/cpu/_02263_ ;
 wire \soc/cpu/_02264_ ;
 wire \soc/cpu/_02265_ ;
 wire \soc/cpu/_02266_ ;
 wire \soc/cpu/_02267_ ;
 wire \soc/cpu/_02268_ ;
 wire \soc/cpu/_02269_ ;
 wire \soc/cpu/_02270_ ;
 wire \soc/cpu/_02271_ ;
 wire \soc/cpu/_02272_ ;
 wire \soc/cpu/_02273_ ;
 wire \soc/cpu/_02274_ ;
 wire \soc/cpu/_02275_ ;
 wire \soc/cpu/_02276_ ;
 wire \soc/cpu/_02277_ ;
 wire \soc/cpu/_02278_ ;
 wire \soc/cpu/_02279_ ;
 wire \soc/cpu/_02280_ ;
 wire \soc/cpu/_02281_ ;
 wire \soc/cpu/_02282_ ;
 wire \soc/cpu/_02283_ ;
 wire \soc/cpu/_02284_ ;
 wire \soc/cpu/_02285_ ;
 wire \soc/cpu/_02286_ ;
 wire \soc/cpu/_02287_ ;
 wire \soc/cpu/_02288_ ;
 wire \soc/cpu/_02289_ ;
 wire \soc/cpu/_02290_ ;
 wire \soc/cpu/_02291_ ;
 wire \soc/cpu/_02292_ ;
 wire \soc/cpu/_02293_ ;
 wire \soc/cpu/_02294_ ;
 wire \soc/cpu/_02295_ ;
 wire net910;
 wire net909;
 wire \soc/cpu/_02298_ ;
 wire \soc/cpu/_02299_ ;
 wire \soc/cpu/_02300_ ;
 wire \soc/cpu/_02301_ ;
 wire \soc/cpu/_02302_ ;
 wire net908;
 wire \soc/cpu/_02304_ ;
 wire net907;
 wire \soc/cpu/_02306_ ;
 wire \soc/cpu/_02307_ ;
 wire \soc/cpu/_02308_ ;
 wire \soc/cpu/_02309_ ;
 wire \soc/cpu/_02310_ ;
 wire \soc/cpu/_02311_ ;
 wire \soc/cpu/_02312_ ;
 wire \soc/cpu/_02313_ ;
 wire net906;
 wire net905;
 wire \soc/cpu/_02316_ ;
 wire \soc/cpu/_02317_ ;
 wire net904;
 wire \soc/cpu/_02319_ ;
 wire \soc/cpu/_02320_ ;
 wire \soc/cpu/_02321_ ;
 wire \soc/cpu/_02322_ ;
 wire \soc/cpu/_02323_ ;
 wire \soc/cpu/_02324_ ;
 wire net903;
 wire \soc/cpu/_02326_ ;
 wire \soc/cpu/_02327_ ;
 wire \soc/cpu/_02328_ ;
 wire \soc/cpu/_02329_ ;
 wire net902;
 wire \soc/cpu/_02331_ ;
 wire \soc/cpu/_02332_ ;
 wire \soc/cpu/_02333_ ;
 wire \soc/cpu/_02334_ ;
 wire \soc/cpu/_02335_ ;
 wire \soc/cpu/_02336_ ;
 wire net901;
 wire \soc/cpu/_02338_ ;
 wire \soc/cpu/_02339_ ;
 wire \soc/cpu/_02340_ ;
 wire \soc/cpu/_02341_ ;
 wire net900;
 wire \soc/cpu/_02343_ ;
 wire \soc/cpu/_02344_ ;
 wire \soc/cpu/_02345_ ;
 wire \soc/cpu/_02346_ ;
 wire \soc/cpu/_02347_ ;
 wire \soc/cpu/_02348_ ;
 wire \soc/cpu/_02349_ ;
 wire \soc/cpu/_02350_ ;
 wire \soc/cpu/_02351_ ;
 wire \soc/cpu/_02352_ ;
 wire \soc/cpu/_02353_ ;
 wire \soc/cpu/_02354_ ;
 wire \soc/cpu/_02355_ ;
 wire \soc/cpu/_02356_ ;
 wire \soc/cpu/_02357_ ;
 wire net899;
 wire net898;
 wire \soc/cpu/_02360_ ;
 wire \soc/cpu/_02361_ ;
 wire \soc/cpu/_02362_ ;
 wire \soc/cpu/_02363_ ;
 wire \soc/cpu/_02364_ ;
 wire \soc/cpu/_02365_ ;
 wire \soc/cpu/_02366_ ;
 wire \soc/cpu/_02367_ ;
 wire net897;
 wire \soc/cpu/_02369_ ;
 wire \soc/cpu/_02370_ ;
 wire \soc/cpu/_02371_ ;
 wire \soc/cpu/_02372_ ;
 wire \soc/cpu/_02373_ ;
 wire \soc/cpu/_02374_ ;
 wire \soc/cpu/_02375_ ;
 wire \soc/cpu/_02376_ ;
 wire \soc/cpu/_02377_ ;
 wire \soc/cpu/_02378_ ;
 wire \soc/cpu/_02379_ ;
 wire \soc/cpu/_02380_ ;
 wire \soc/cpu/_02381_ ;
 wire \soc/cpu/_02382_ ;
 wire net896;
 wire \soc/cpu/_02384_ ;
 wire net895;
 wire \soc/cpu/_02386_ ;
 wire \soc/cpu/_02387_ ;
 wire \soc/cpu/_02388_ ;
 wire \soc/cpu/_02389_ ;
 wire \soc/cpu/_02390_ ;
 wire net894;
 wire \soc/cpu/_02392_ ;
 wire \soc/cpu/_02393_ ;
 wire \soc/cpu/_02394_ ;
 wire \soc/cpu/_02395_ ;
 wire \soc/cpu/_02396_ ;
 wire \soc/cpu/_02397_ ;
 wire \soc/cpu/_02398_ ;
 wire \soc/cpu/_02399_ ;
 wire \soc/cpu/_02400_ ;
 wire \soc/cpu/_02401_ ;
 wire \soc/cpu/_02402_ ;
 wire \soc/cpu/_02403_ ;
 wire \soc/cpu/_02404_ ;
 wire \soc/cpu/_02405_ ;
 wire \soc/cpu/_02406_ ;
 wire \soc/cpu/_02407_ ;
 wire \soc/cpu/_02408_ ;
 wire net893;
 wire net892;
 wire \soc/cpu/_02411_ ;
 wire \soc/cpu/_02412_ ;
 wire net891;
 wire net890;
 wire \soc/cpu/_02415_ ;
 wire \soc/cpu/_02416_ ;
 wire \soc/cpu/_02417_ ;
 wire \soc/cpu/_02418_ ;
 wire \soc/cpu/_02419_ ;
 wire \soc/cpu/_02420_ ;
 wire \soc/cpu/_02421_ ;
 wire \soc/cpu/_02422_ ;
 wire \soc/cpu/_02423_ ;
 wire \soc/cpu/_02424_ ;
 wire \soc/cpu/_02425_ ;
 wire \soc/cpu/_02426_ ;
 wire \soc/cpu/_02427_ ;
 wire \soc/cpu/_02428_ ;
 wire \soc/cpu/_02429_ ;
 wire \soc/cpu/_02430_ ;
 wire \soc/cpu/_02431_ ;
 wire net889;
 wire net888;
 wire net887;
 wire \soc/cpu/_02435_ ;
 wire \soc/cpu/_02436_ ;
 wire \soc/cpu/_02437_ ;
 wire \soc/cpu/_02438_ ;
 wire \soc/cpu/_02439_ ;
 wire \soc/cpu/_02440_ ;
 wire \soc/cpu/_02441_ ;
 wire net886;
 wire \soc/cpu/_02443_ ;
 wire \soc/cpu/_02444_ ;
 wire \soc/cpu/_02445_ ;
 wire \soc/cpu/_02446_ ;
 wire net885;
 wire \soc/cpu/_02448_ ;
 wire \soc/cpu/_02449_ ;
 wire \soc/cpu/_02450_ ;
 wire net884;
 wire \soc/cpu/_02452_ ;
 wire \soc/cpu/_02453_ ;
 wire \soc/cpu/_02454_ ;
 wire net883;
 wire \soc/cpu/_02456_ ;
 wire \soc/cpu/_02457_ ;
 wire \soc/cpu/_02458_ ;
 wire \soc/cpu/_02459_ ;
 wire net882;
 wire \soc/cpu/_02461_ ;
 wire \soc/cpu/_02462_ ;
 wire \soc/cpu/_02463_ ;
 wire \soc/cpu/_02464_ ;
 wire \soc/cpu/_02465_ ;
 wire \soc/cpu/_02466_ ;
 wire \soc/cpu/_02467_ ;
 wire \soc/cpu/_02468_ ;
 wire \soc/cpu/_02469_ ;
 wire \soc/cpu/_02470_ ;
 wire \soc/cpu/_02471_ ;
 wire net881;
 wire \soc/cpu/_02473_ ;
 wire \soc/cpu/_02474_ ;
 wire \soc/cpu/_02475_ ;
 wire \soc/cpu/_02476_ ;
 wire \soc/cpu/_02477_ ;
 wire \soc/cpu/_02478_ ;
 wire \soc/cpu/_02479_ ;
 wire \soc/cpu/_02480_ ;
 wire \soc/cpu/_02481_ ;
 wire \soc/cpu/_02482_ ;
 wire \soc/cpu/_02483_ ;
 wire \soc/cpu/_02484_ ;
 wire \soc/cpu/_02485_ ;
 wire \soc/cpu/_02486_ ;
 wire \soc/cpu/_02487_ ;
 wire \soc/cpu/_02488_ ;
 wire \soc/cpu/_02489_ ;
 wire \soc/cpu/_02490_ ;
 wire \soc/cpu/_02491_ ;
 wire \soc/cpu/_02492_ ;
 wire \soc/cpu/_02493_ ;
 wire \soc/cpu/_02494_ ;
 wire \soc/cpu/_02495_ ;
 wire \soc/cpu/_02496_ ;
 wire \soc/cpu/_02497_ ;
 wire \soc/cpu/_02498_ ;
 wire net880;
 wire \soc/cpu/_02500_ ;
 wire \soc/cpu/_02501_ ;
 wire net879;
 wire \soc/cpu/_02503_ ;
 wire \soc/cpu/_02504_ ;
 wire \soc/cpu/_02505_ ;
 wire \soc/cpu/_02506_ ;
 wire \soc/cpu/_02507_ ;
 wire \soc/cpu/_02508_ ;
 wire \soc/cpu/_02509_ ;
 wire net878;
 wire \soc/cpu/_02511_ ;
 wire net877;
 wire \soc/cpu/_02513_ ;
 wire \soc/cpu/_02514_ ;
 wire \soc/cpu/_02515_ ;
 wire \soc/cpu/_02516_ ;
 wire \soc/cpu/_02517_ ;
 wire \soc/cpu/_02518_ ;
 wire \soc/cpu/_02519_ ;
 wire \soc/cpu/_02520_ ;
 wire \soc/cpu/_02521_ ;
 wire net876;
 wire \soc/cpu/_02523_ ;
 wire \soc/cpu/_02524_ ;
 wire \soc/cpu/_02525_ ;
 wire \soc/cpu/_02526_ ;
 wire \soc/cpu/_02527_ ;
 wire \soc/cpu/_02528_ ;
 wire \soc/cpu/_02529_ ;
 wire \soc/cpu/_02530_ ;
 wire \soc/cpu/_02531_ ;
 wire \soc/cpu/_02532_ ;
 wire net875;
 wire net874;
 wire \soc/cpu/_02535_ ;
 wire \soc/cpu/_02536_ ;
 wire \soc/cpu/_02537_ ;
 wire \soc/cpu/_02538_ ;
 wire net873;
 wire \soc/cpu/_02540_ ;
 wire net872;
 wire \soc/cpu/_02542_ ;
 wire net871;
 wire \soc/cpu/_02544_ ;
 wire net870;
 wire \soc/cpu/_02546_ ;
 wire \soc/cpu/_02547_ ;
 wire \soc/cpu/_02548_ ;
 wire \soc/cpu/_02549_ ;
 wire \soc/cpu/_02550_ ;
 wire net869;
 wire \soc/cpu/_02552_ ;
 wire \soc/cpu/_02553_ ;
 wire \soc/cpu/_02554_ ;
 wire net868;
 wire net867;
 wire \soc/cpu/_02557_ ;
 wire \soc/cpu/_02558_ ;
 wire net866;
 wire \soc/cpu/_02560_ ;
 wire \soc/cpu/_02561_ ;
 wire \soc/cpu/_02562_ ;
 wire \soc/cpu/_02563_ ;
 wire \soc/cpu/_02564_ ;
 wire \soc/cpu/_02565_ ;
 wire \soc/cpu/_02566_ ;
 wire net865;
 wire \soc/cpu/_02568_ ;
 wire \soc/cpu/_02569_ ;
 wire \soc/cpu/_02570_ ;
 wire \soc/cpu/_02571_ ;
 wire \soc/cpu/_02572_ ;
 wire \soc/cpu/_02573_ ;
 wire \soc/cpu/_02574_ ;
 wire \soc/cpu/_02575_ ;
 wire \soc/cpu/_02576_ ;
 wire \soc/cpu/_02577_ ;
 wire \soc/cpu/_02578_ ;
 wire \soc/cpu/_02579_ ;
 wire \soc/cpu/_02580_ ;
 wire \soc/cpu/_02581_ ;
 wire \soc/cpu/_02582_ ;
 wire \soc/cpu/_02583_ ;
 wire \soc/cpu/_02584_ ;
 wire \soc/cpu/_02585_ ;
 wire \soc/cpu/_02586_ ;
 wire \soc/cpu/_02587_ ;
 wire \soc/cpu/_02588_ ;
 wire \soc/cpu/_02589_ ;
 wire \soc/cpu/_02590_ ;
 wire \soc/cpu/_02591_ ;
 wire \soc/cpu/_02592_ ;
 wire \soc/cpu/_02593_ ;
 wire \soc/cpu/_02594_ ;
 wire \soc/cpu/_02595_ ;
 wire \soc/cpu/_02596_ ;
 wire \soc/cpu/_02597_ ;
 wire \soc/cpu/_02598_ ;
 wire \soc/cpu/_02599_ ;
 wire \soc/cpu/_02600_ ;
 wire \soc/cpu/_02601_ ;
 wire \soc/cpu/_02602_ ;
 wire \soc/cpu/_02603_ ;
 wire \soc/cpu/_02604_ ;
 wire \soc/cpu/_02605_ ;
 wire \soc/cpu/_02606_ ;
 wire net864;
 wire \soc/cpu/_02608_ ;
 wire \soc/cpu/_02609_ ;
 wire \soc/cpu/_02610_ ;
 wire \soc/cpu/_02611_ ;
 wire \soc/cpu/_02612_ ;
 wire \soc/cpu/_02613_ ;
 wire \soc/cpu/_02614_ ;
 wire \soc/cpu/_02615_ ;
 wire \soc/cpu/_02616_ ;
 wire \soc/cpu/_02617_ ;
 wire \soc/cpu/_02618_ ;
 wire \soc/cpu/_02619_ ;
 wire \soc/cpu/_02620_ ;
 wire \soc/cpu/_02621_ ;
 wire \soc/cpu/_02622_ ;
 wire \soc/cpu/_02623_ ;
 wire \soc/cpu/_02624_ ;
 wire \soc/cpu/_02625_ ;
 wire \soc/cpu/_02626_ ;
 wire \soc/cpu/_02627_ ;
 wire \soc/cpu/_02628_ ;
 wire \soc/cpu/_02629_ ;
 wire \soc/cpu/_02630_ ;
 wire \soc/cpu/_02631_ ;
 wire \soc/cpu/_02632_ ;
 wire \soc/cpu/_02633_ ;
 wire \soc/cpu/_02634_ ;
 wire \soc/cpu/_02635_ ;
 wire \soc/cpu/_02636_ ;
 wire \soc/cpu/_02637_ ;
 wire \soc/cpu/_02638_ ;
 wire \soc/cpu/_02639_ ;
 wire \soc/cpu/_02640_ ;
 wire \soc/cpu/_02641_ ;
 wire \soc/cpu/_02642_ ;
 wire \soc/cpu/_02643_ ;
 wire \soc/cpu/_02644_ ;
 wire \soc/cpu/_02645_ ;
 wire \soc/cpu/_02646_ ;
 wire \soc/cpu/_02647_ ;
 wire \soc/cpu/_02648_ ;
 wire \soc/cpu/_02649_ ;
 wire \soc/cpu/_02650_ ;
 wire \soc/cpu/_02651_ ;
 wire \soc/cpu/_02652_ ;
 wire \soc/cpu/_02653_ ;
 wire \soc/cpu/_02654_ ;
 wire \soc/cpu/_02655_ ;
 wire \soc/cpu/_02656_ ;
 wire \soc/cpu/_02657_ ;
 wire \soc/cpu/_02658_ ;
 wire \soc/cpu/_02659_ ;
 wire \soc/cpu/_02660_ ;
 wire \soc/cpu/_02661_ ;
 wire \soc/cpu/_02662_ ;
 wire \soc/cpu/_02663_ ;
 wire \soc/cpu/_02664_ ;
 wire \soc/cpu/_02665_ ;
 wire \soc/cpu/_02666_ ;
 wire \soc/cpu/_02667_ ;
 wire \soc/cpu/_02668_ ;
 wire \soc/cpu/_02669_ ;
 wire \soc/cpu/_02670_ ;
 wire \soc/cpu/_02671_ ;
 wire \soc/cpu/_02672_ ;
 wire \soc/cpu/_02673_ ;
 wire \soc/cpu/_02674_ ;
 wire \soc/cpu/_02675_ ;
 wire \soc/cpu/_02676_ ;
 wire \soc/cpu/_02677_ ;
 wire \soc/cpu/_02678_ ;
 wire \soc/cpu/_02679_ ;
 wire \soc/cpu/_02680_ ;
 wire \soc/cpu/_02681_ ;
 wire \soc/cpu/_02682_ ;
 wire \soc/cpu/_02683_ ;
 wire \soc/cpu/_02684_ ;
 wire \soc/cpu/_02685_ ;
 wire \soc/cpu/_02686_ ;
 wire \soc/cpu/_02687_ ;
 wire \soc/cpu/_02688_ ;
 wire \soc/cpu/_02689_ ;
 wire \soc/cpu/_02690_ ;
 wire \soc/cpu/_02691_ ;
 wire \soc/cpu/_02692_ ;
 wire net863;
 wire \soc/cpu/_02694_ ;
 wire \soc/cpu/_02695_ ;
 wire \soc/cpu/_02696_ ;
 wire net862;
 wire \soc/cpu/_02698_ ;
 wire \soc/cpu/_02699_ ;
 wire net861;
 wire \soc/cpu/_02701_ ;
 wire \soc/cpu/_02702_ ;
 wire net860;
 wire \soc/cpu/_02704_ ;
 wire \soc/cpu/_02705_ ;
 wire net859;
 wire \soc/cpu/_02707_ ;
 wire \soc/cpu/_02708_ ;
 wire \soc/cpu/_02709_ ;
 wire \soc/cpu/_02710_ ;
 wire \soc/cpu/_02711_ ;
 wire \soc/cpu/_02712_ ;
 wire net858;
 wire net857;
 wire net856;
 wire \soc/cpu/_02716_ ;
 wire \soc/cpu/_02717_ ;
 wire \soc/cpu/_02718_ ;
 wire \soc/cpu/_02719_ ;
 wire \soc/cpu/_02720_ ;
 wire \soc/cpu/_02721_ ;
 wire \soc/cpu/_02722_ ;
 wire \soc/cpu/_02723_ ;
 wire \soc/cpu/_02724_ ;
 wire \soc/cpu/_02725_ ;
 wire \soc/cpu/_02726_ ;
 wire \soc/cpu/_02727_ ;
 wire \soc/cpu/_02728_ ;
 wire \soc/cpu/_02729_ ;
 wire \soc/cpu/_02730_ ;
 wire \soc/cpu/_02731_ ;
 wire \soc/cpu/_02732_ ;
 wire \soc/cpu/_02733_ ;
 wire \soc/cpu/_02734_ ;
 wire \soc/cpu/_02735_ ;
 wire \soc/cpu/_02736_ ;
 wire \soc/cpu/_02737_ ;
 wire \soc/cpu/_02738_ ;
 wire \soc/cpu/_02739_ ;
 wire \soc/cpu/_02740_ ;
 wire \soc/cpu/_02741_ ;
 wire \soc/cpu/_02742_ ;
 wire \soc/cpu/_02743_ ;
 wire \soc/cpu/_02744_ ;
 wire \soc/cpu/_02745_ ;
 wire \soc/cpu/_02746_ ;
 wire \soc/cpu/_02747_ ;
 wire \soc/cpu/_02748_ ;
 wire \soc/cpu/_02749_ ;
 wire \soc/cpu/_02750_ ;
 wire \soc/cpu/_02751_ ;
 wire \soc/cpu/_02752_ ;
 wire \soc/cpu/_02753_ ;
 wire \soc/cpu/_02754_ ;
 wire \soc/cpu/_02755_ ;
 wire \soc/cpu/_02756_ ;
 wire \soc/cpu/_02757_ ;
 wire \soc/cpu/_02758_ ;
 wire \soc/cpu/_02759_ ;
 wire \soc/cpu/_02760_ ;
 wire \soc/cpu/_02761_ ;
 wire \soc/cpu/_02762_ ;
 wire \soc/cpu/_02763_ ;
 wire \soc/cpu/_02764_ ;
 wire net855;
 wire \soc/cpu/_02766_ ;
 wire net854;
 wire \soc/cpu/_02768_ ;
 wire net853;
 wire net852;
 wire \soc/cpu/_02771_ ;
 wire \soc/cpu/_02772_ ;
 wire \soc/cpu/_02773_ ;
 wire \soc/cpu/_02774_ ;
 wire \soc/cpu/_02775_ ;
 wire \soc/cpu/_02776_ ;
 wire \soc/cpu/_02777_ ;
 wire \soc/cpu/_02778_ ;
 wire \soc/cpu/_02779_ ;
 wire \soc/cpu/_02780_ ;
 wire net851;
 wire \soc/cpu/_02782_ ;
 wire \soc/cpu/_02783_ ;
 wire \soc/cpu/_02784_ ;
 wire \soc/cpu/_02785_ ;
 wire \soc/cpu/_02786_ ;
 wire \soc/cpu/_02787_ ;
 wire \soc/cpu/_02788_ ;
 wire \soc/cpu/_02789_ ;
 wire \soc/cpu/_02790_ ;
 wire \soc/cpu/_02791_ ;
 wire \soc/cpu/_02792_ ;
 wire \soc/cpu/_02793_ ;
 wire \soc/cpu/_02794_ ;
 wire \soc/cpu/_02795_ ;
 wire \soc/cpu/_02796_ ;
 wire net850;
 wire \soc/cpu/_02798_ ;
 wire \soc/cpu/_02799_ ;
 wire net849;
 wire \soc/cpu/_02801_ ;
 wire \soc/cpu/_02802_ ;
 wire \soc/cpu/_02803_ ;
 wire \soc/cpu/_02804_ ;
 wire \soc/cpu/_02805_ ;
 wire \soc/cpu/_02806_ ;
 wire \soc/cpu/_02807_ ;
 wire \soc/cpu/_02808_ ;
 wire \soc/cpu/_02809_ ;
 wire \soc/cpu/_02810_ ;
 wire \soc/cpu/_02811_ ;
 wire \soc/cpu/_02812_ ;
 wire \soc/cpu/_02813_ ;
 wire net848;
 wire \soc/cpu/_02815_ ;
 wire \soc/cpu/_02816_ ;
 wire \soc/cpu/_02817_ ;
 wire net847;
 wire \soc/cpu/_02819_ ;
 wire net846;
 wire net845;
 wire \soc/cpu/_02822_ ;
 wire \soc/cpu/_02823_ ;
 wire net844;
 wire \soc/cpu/_02825_ ;
 wire \soc/cpu/_02826_ ;
 wire \soc/cpu/_02827_ ;
 wire \soc/cpu/_02828_ ;
 wire \soc/cpu/_02829_ ;
 wire \soc/cpu/_02830_ ;
 wire \soc/cpu/_02831_ ;
 wire \soc/cpu/_02832_ ;
 wire \soc/cpu/_02833_ ;
 wire \soc/cpu/_02834_ ;
 wire \soc/cpu/_02835_ ;
 wire \soc/cpu/_02836_ ;
 wire \soc/cpu/_02837_ ;
 wire \soc/cpu/_02838_ ;
 wire \soc/cpu/_02839_ ;
 wire \soc/cpu/_02840_ ;
 wire \soc/cpu/_02841_ ;
 wire \soc/cpu/_02842_ ;
 wire \soc/cpu/_02843_ ;
 wire \soc/cpu/_02844_ ;
 wire \soc/cpu/_02845_ ;
 wire \soc/cpu/_02846_ ;
 wire \soc/cpu/_02847_ ;
 wire \soc/cpu/_02848_ ;
 wire \soc/cpu/_02849_ ;
 wire \soc/cpu/_02850_ ;
 wire \soc/cpu/_02851_ ;
 wire \soc/cpu/_02852_ ;
 wire \soc/cpu/_02853_ ;
 wire net843;
 wire \soc/cpu/_02855_ ;
 wire \soc/cpu/_02856_ ;
 wire \soc/cpu/_02857_ ;
 wire net842;
 wire \soc/cpu/_02859_ ;
 wire \soc/cpu/_02860_ ;
 wire \soc/cpu/_02861_ ;
 wire \soc/cpu/_02862_ ;
 wire \soc/cpu/_02863_ ;
 wire \soc/cpu/_02864_ ;
 wire \soc/cpu/_02865_ ;
 wire \soc/cpu/_02866_ ;
 wire \soc/cpu/_02867_ ;
 wire \soc/cpu/_02868_ ;
 wire \soc/cpu/_02869_ ;
 wire \soc/cpu/_02870_ ;
 wire \soc/cpu/_02871_ ;
 wire \soc/cpu/_02872_ ;
 wire \soc/cpu/_02873_ ;
 wire \soc/cpu/_02874_ ;
 wire \soc/cpu/_02875_ ;
 wire \soc/cpu/_02876_ ;
 wire \soc/cpu/_02877_ ;
 wire \soc/cpu/_02878_ ;
 wire \soc/cpu/_02879_ ;
 wire \soc/cpu/_02880_ ;
 wire \soc/cpu/_02881_ ;
 wire \soc/cpu/_02882_ ;
 wire net841;
 wire \soc/cpu/_02884_ ;
 wire \soc/cpu/_02885_ ;
 wire \soc/cpu/_02886_ ;
 wire \soc/cpu/_02887_ ;
 wire \soc/cpu/_02888_ ;
 wire \soc/cpu/_02889_ ;
 wire net840;
 wire net839;
 wire \soc/cpu/_02892_ ;
 wire \soc/cpu/_02893_ ;
 wire \soc/cpu/_02894_ ;
 wire \soc/cpu/_02895_ ;
 wire \soc/cpu/_02896_ ;
 wire \soc/cpu/_02897_ ;
 wire \soc/cpu/_02898_ ;
 wire \soc/cpu/_02899_ ;
 wire net838;
 wire \soc/cpu/_02901_ ;
 wire \soc/cpu/_02902_ ;
 wire \soc/cpu/_02903_ ;
 wire \soc/cpu/_02904_ ;
 wire net837;
 wire \soc/cpu/_02906_ ;
 wire net836;
 wire net835;
 wire \soc/cpu/_02909_ ;
 wire \soc/cpu/_02910_ ;
 wire \soc/cpu/_02911_ ;
 wire net834;
 wire net833;
 wire net832;
 wire net831;
 wire \soc/cpu/_02916_ ;
 wire \soc/cpu/_02917_ ;
 wire \soc/cpu/_02918_ ;
 wire \soc/cpu/_02919_ ;
 wire \soc/cpu/_02920_ ;
 wire \soc/cpu/_02921_ ;
 wire \soc/cpu/_02922_ ;
 wire net830;
 wire \soc/cpu/_02924_ ;
 wire \soc/cpu/_02925_ ;
 wire \soc/cpu/_02926_ ;
 wire \soc/cpu/_02927_ ;
 wire net829;
 wire \soc/cpu/_02929_ ;
 wire \soc/cpu/_02930_ ;
 wire \soc/cpu/_02931_ ;
 wire net828;
 wire net827;
 wire net826;
 wire \soc/cpu/_02935_ ;
 wire net825;
 wire \soc/cpu/_02937_ ;
 wire \soc/cpu/_02938_ ;
 wire net824;
 wire \soc/cpu/_02940_ ;
 wire net823;
 wire \soc/cpu/_02942_ ;
 wire net822;
 wire \soc/cpu/_02944_ ;
 wire \soc/cpu/_02945_ ;
 wire \soc/cpu/_02946_ ;
 wire \soc/cpu/_02947_ ;
 wire net821;
 wire \soc/cpu/_02949_ ;
 wire \soc/cpu/_02950_ ;
 wire \soc/cpu/_02951_ ;
 wire \soc/cpu/_02952_ ;
 wire \soc/cpu/_02953_ ;
 wire \soc/cpu/_02954_ ;
 wire \soc/cpu/_02955_ ;
 wire net820;
 wire \soc/cpu/_02957_ ;
 wire \soc/cpu/_02958_ ;
 wire \soc/cpu/_02959_ ;
 wire \soc/cpu/_02960_ ;
 wire \soc/cpu/_02961_ ;
 wire \soc/cpu/_02962_ ;
 wire \soc/cpu/_02963_ ;
 wire \soc/cpu/_02964_ ;
 wire \soc/cpu/_02965_ ;
 wire \soc/cpu/_02966_ ;
 wire \soc/cpu/_02967_ ;
 wire \soc/cpu/_02968_ ;
 wire \soc/cpu/_02969_ ;
 wire \soc/cpu/_02970_ ;
 wire \soc/cpu/_02971_ ;
 wire \soc/cpu/_02972_ ;
 wire \soc/cpu/_02973_ ;
 wire net819;
 wire \soc/cpu/_02975_ ;
 wire \soc/cpu/_02976_ ;
 wire net818;
 wire \soc/cpu/_02978_ ;
 wire \soc/cpu/_02979_ ;
 wire \soc/cpu/_02980_ ;
 wire \soc/cpu/_02981_ ;
 wire \soc/cpu/_02982_ ;
 wire \soc/cpu/_02983_ ;
 wire \soc/cpu/_02984_ ;
 wire \soc/cpu/_02985_ ;
 wire net817;
 wire \soc/cpu/_02987_ ;
 wire \soc/cpu/_02988_ ;
 wire \soc/cpu/_02989_ ;
 wire net816;
 wire \soc/cpu/_02991_ ;
 wire \soc/cpu/_02992_ ;
 wire \soc/cpu/_02993_ ;
 wire \soc/cpu/_02994_ ;
 wire \soc/cpu/_02995_ ;
 wire \soc/cpu/_02996_ ;
 wire \soc/cpu/_02997_ ;
 wire \soc/cpu/_02998_ ;
 wire \soc/cpu/_02999_ ;
 wire \soc/cpu/_03000_ ;
 wire \soc/cpu/_03001_ ;
 wire \soc/cpu/_03002_ ;
 wire \soc/cpu/_03003_ ;
 wire \soc/cpu/_03004_ ;
 wire \soc/cpu/_03005_ ;
 wire \soc/cpu/_03006_ ;
 wire \soc/cpu/_03007_ ;
 wire \soc/cpu/_03008_ ;
 wire \soc/cpu/_03009_ ;
 wire \soc/cpu/_03010_ ;
 wire \soc/cpu/_03011_ ;
 wire \soc/cpu/_03012_ ;
 wire \soc/cpu/_03013_ ;
 wire \soc/cpu/_03014_ ;
 wire \soc/cpu/_03015_ ;
 wire \soc/cpu/_03016_ ;
 wire \soc/cpu/_03017_ ;
 wire \soc/cpu/_03018_ ;
 wire \soc/cpu/_03019_ ;
 wire net815;
 wire \soc/cpu/_03021_ ;
 wire \soc/cpu/_03022_ ;
 wire \soc/cpu/_03023_ ;
 wire \soc/cpu/_03024_ ;
 wire \soc/cpu/_03025_ ;
 wire \soc/cpu/_03026_ ;
 wire \soc/cpu/_03027_ ;
 wire \soc/cpu/_03028_ ;
 wire \soc/cpu/_03029_ ;
 wire \soc/cpu/_03030_ ;
 wire \soc/cpu/_03031_ ;
 wire \soc/cpu/_03032_ ;
 wire \soc/cpu/_03033_ ;
 wire \soc/cpu/_03034_ ;
 wire \soc/cpu/_03035_ ;
 wire \soc/cpu/_03036_ ;
 wire \soc/cpu/_03037_ ;
 wire \soc/cpu/_03038_ ;
 wire \soc/cpu/_03039_ ;
 wire \soc/cpu/_03040_ ;
 wire \soc/cpu/_03041_ ;
 wire \soc/cpu/_03042_ ;
 wire \soc/cpu/_03043_ ;
 wire \soc/cpu/_03044_ ;
 wire \soc/cpu/_03045_ ;
 wire \soc/cpu/_03046_ ;
 wire \soc/cpu/_03047_ ;
 wire \soc/cpu/_03048_ ;
 wire \soc/cpu/_03049_ ;
 wire \soc/cpu/_03050_ ;
 wire \soc/cpu/_03051_ ;
 wire \soc/cpu/_03052_ ;
 wire \soc/cpu/_03053_ ;
 wire \soc/cpu/_03054_ ;
 wire \soc/cpu/_03055_ ;
 wire \soc/cpu/_03056_ ;
 wire \soc/cpu/_03057_ ;
 wire \soc/cpu/_03058_ ;
 wire \soc/cpu/_03059_ ;
 wire \soc/cpu/_03060_ ;
 wire \soc/cpu/_03061_ ;
 wire \soc/cpu/_03062_ ;
 wire \soc/cpu/_03063_ ;
 wire \soc/cpu/_03064_ ;
 wire \soc/cpu/_03065_ ;
 wire \soc/cpu/_03066_ ;
 wire \soc/cpu/_03067_ ;
 wire \soc/cpu/_03068_ ;
 wire \soc/cpu/_03069_ ;
 wire \soc/cpu/_03070_ ;
 wire \soc/cpu/_03071_ ;
 wire \soc/cpu/_03072_ ;
 wire \soc/cpu/_03073_ ;
 wire \soc/cpu/_03074_ ;
 wire \soc/cpu/_03075_ ;
 wire \soc/cpu/_03076_ ;
 wire \soc/cpu/_03077_ ;
 wire \soc/cpu/_03078_ ;
 wire \soc/cpu/_03079_ ;
 wire \soc/cpu/_03080_ ;
 wire \soc/cpu/_03081_ ;
 wire \soc/cpu/_03082_ ;
 wire \soc/cpu/_03083_ ;
 wire \soc/cpu/_03084_ ;
 wire \soc/cpu/_03085_ ;
 wire \soc/cpu/_03086_ ;
 wire \soc/cpu/_03087_ ;
 wire \soc/cpu/_03088_ ;
 wire \soc/cpu/_03089_ ;
 wire \soc/cpu/_03090_ ;
 wire \soc/cpu/_03091_ ;
 wire \soc/cpu/_03092_ ;
 wire \soc/cpu/_03093_ ;
 wire \soc/cpu/_03094_ ;
 wire \soc/cpu/_03095_ ;
 wire \soc/cpu/_03096_ ;
 wire \soc/cpu/_03097_ ;
 wire \soc/cpu/_03098_ ;
 wire \soc/cpu/_03099_ ;
 wire \soc/cpu/_03100_ ;
 wire \soc/cpu/_03101_ ;
 wire \soc/cpu/_03102_ ;
 wire \soc/cpu/_03103_ ;
 wire \soc/cpu/_03104_ ;
 wire \soc/cpu/_03105_ ;
 wire \soc/cpu/_03106_ ;
 wire \soc/cpu/_03107_ ;
 wire \soc/cpu/_03108_ ;
 wire \soc/cpu/_03109_ ;
 wire \soc/cpu/_03110_ ;
 wire \soc/cpu/_03111_ ;
 wire \soc/cpu/_03112_ ;
 wire \soc/cpu/_03113_ ;
 wire \soc/cpu/_03114_ ;
 wire \soc/cpu/_03115_ ;
 wire \soc/cpu/_03116_ ;
 wire \soc/cpu/_03117_ ;
 wire \soc/cpu/_03118_ ;
 wire \soc/cpu/_03119_ ;
 wire \soc/cpu/_03120_ ;
 wire \soc/cpu/_03121_ ;
 wire \soc/cpu/_03122_ ;
 wire \soc/cpu/_03123_ ;
 wire \soc/cpu/_03124_ ;
 wire \soc/cpu/_03125_ ;
 wire \soc/cpu/_03126_ ;
 wire \soc/cpu/_03127_ ;
 wire \soc/cpu/_03128_ ;
 wire \soc/cpu/_03129_ ;
 wire \soc/cpu/_03130_ ;
 wire \soc/cpu/_03131_ ;
 wire \soc/cpu/_03132_ ;
 wire \soc/cpu/_03133_ ;
 wire \soc/cpu/_03134_ ;
 wire net814;
 wire \soc/cpu/_03136_ ;
 wire \soc/cpu/_03137_ ;
 wire \soc/cpu/_03138_ ;
 wire \soc/cpu/_03139_ ;
 wire \soc/cpu/_03140_ ;
 wire \soc/cpu/_03141_ ;
 wire \soc/cpu/_03142_ ;
 wire \soc/cpu/_03143_ ;
 wire \soc/cpu/_03144_ ;
 wire \soc/cpu/_03145_ ;
 wire \soc/cpu/_03146_ ;
 wire \soc/cpu/_03147_ ;
 wire \soc/cpu/_03148_ ;
 wire \soc/cpu/_03149_ ;
 wire \soc/cpu/_03150_ ;
 wire \soc/cpu/_03151_ ;
 wire \soc/cpu/_03152_ ;
 wire \soc/cpu/_03153_ ;
 wire \soc/cpu/_03154_ ;
 wire \soc/cpu/_03155_ ;
 wire \soc/cpu/_03156_ ;
 wire \soc/cpu/_03157_ ;
 wire \soc/cpu/_03158_ ;
 wire \soc/cpu/_03159_ ;
 wire \soc/cpu/_03160_ ;
 wire \soc/cpu/_03161_ ;
 wire \soc/cpu/_03162_ ;
 wire \soc/cpu/_03163_ ;
 wire \soc/cpu/_03164_ ;
 wire \soc/cpu/_03165_ ;
 wire \soc/cpu/_03166_ ;
 wire \soc/cpu/_03167_ ;
 wire \soc/cpu/_03168_ ;
 wire \soc/cpu/_03169_ ;
 wire \soc/cpu/_03170_ ;
 wire \soc/cpu/_03171_ ;
 wire \soc/cpu/_03172_ ;
 wire \soc/cpu/_03173_ ;
 wire \soc/cpu/_03174_ ;
 wire \soc/cpu/_03175_ ;
 wire \soc/cpu/_03176_ ;
 wire \soc/cpu/_03177_ ;
 wire \soc/cpu/_03178_ ;
 wire \soc/cpu/_03179_ ;
 wire \soc/cpu/_03180_ ;
 wire \soc/cpu/_03181_ ;
 wire \soc/cpu/_03182_ ;
 wire \soc/cpu/_03183_ ;
 wire \soc/cpu/_03184_ ;
 wire \soc/cpu/_03185_ ;
 wire \soc/cpu/_03186_ ;
 wire \soc/cpu/_03187_ ;
 wire \soc/cpu/_03188_ ;
 wire \soc/cpu/_03189_ ;
 wire \soc/cpu/_03190_ ;
 wire \soc/cpu/_03191_ ;
 wire \soc/cpu/_03192_ ;
 wire \soc/cpu/_03193_ ;
 wire \soc/cpu/_03194_ ;
 wire \soc/cpu/_03195_ ;
 wire \soc/cpu/_03196_ ;
 wire \soc/cpu/_03197_ ;
 wire \soc/cpu/_03198_ ;
 wire \soc/cpu/_03199_ ;
 wire \soc/cpu/_03200_ ;
 wire \soc/cpu/_03201_ ;
 wire \soc/cpu/_03202_ ;
 wire \soc/cpu/_03203_ ;
 wire \soc/cpu/_03204_ ;
 wire \soc/cpu/_03205_ ;
 wire \soc/cpu/_03206_ ;
 wire \soc/cpu/_03207_ ;
 wire \soc/cpu/_03208_ ;
 wire \soc/cpu/_03209_ ;
 wire \soc/cpu/_03210_ ;
 wire \soc/cpu/_03211_ ;
 wire \soc/cpu/_03212_ ;
 wire \soc/cpu/_03213_ ;
 wire \soc/cpu/_03214_ ;
 wire \soc/cpu/_03215_ ;
 wire \soc/cpu/_03216_ ;
 wire \soc/cpu/_03217_ ;
 wire \soc/cpu/_03218_ ;
 wire \soc/cpu/_03219_ ;
 wire \soc/cpu/_03220_ ;
 wire \soc/cpu/_03221_ ;
 wire \soc/cpu/_03222_ ;
 wire \soc/cpu/_03223_ ;
 wire \soc/cpu/_03224_ ;
 wire \soc/cpu/_03225_ ;
 wire \soc/cpu/_03226_ ;
 wire \soc/cpu/_03227_ ;
 wire \soc/cpu/_03228_ ;
 wire \soc/cpu/_03229_ ;
 wire \soc/cpu/_03230_ ;
 wire \soc/cpu/_03231_ ;
 wire \soc/cpu/_03232_ ;
 wire \soc/cpu/_03233_ ;
 wire \soc/cpu/_03234_ ;
 wire \soc/cpu/_03235_ ;
 wire \soc/cpu/_03236_ ;
 wire \soc/cpu/_03237_ ;
 wire \soc/cpu/_03238_ ;
 wire \soc/cpu/_03239_ ;
 wire \soc/cpu/_03240_ ;
 wire \soc/cpu/_03241_ ;
 wire \soc/cpu/_03242_ ;
 wire \soc/cpu/_03243_ ;
 wire \soc/cpu/_03244_ ;
 wire \soc/cpu/_03245_ ;
 wire \soc/cpu/_03246_ ;
 wire \soc/cpu/_03247_ ;
 wire \soc/cpu/_03248_ ;
 wire \soc/cpu/_03249_ ;
 wire \soc/cpu/_03250_ ;
 wire \soc/cpu/_03251_ ;
 wire \soc/cpu/_03252_ ;
 wire \soc/cpu/_03253_ ;
 wire \soc/cpu/_03254_ ;
 wire \soc/cpu/_03255_ ;
 wire \soc/cpu/_03256_ ;
 wire \soc/cpu/_03257_ ;
 wire \soc/cpu/_03258_ ;
 wire \soc/cpu/_03259_ ;
 wire \soc/cpu/_03260_ ;
 wire \soc/cpu/_03261_ ;
 wire \soc/cpu/_03262_ ;
 wire \soc/cpu/_03263_ ;
 wire \soc/cpu/_03264_ ;
 wire \soc/cpu/_03265_ ;
 wire \soc/cpu/_03266_ ;
 wire \soc/cpu/_03267_ ;
 wire \soc/cpu/_03268_ ;
 wire \soc/cpu/_03269_ ;
 wire \soc/cpu/_03270_ ;
 wire \soc/cpu/_03271_ ;
 wire \soc/cpu/_03272_ ;
 wire \soc/cpu/_03273_ ;
 wire \soc/cpu/_03274_ ;
 wire \soc/cpu/_03275_ ;
 wire \soc/cpu/_03276_ ;
 wire \soc/cpu/_03277_ ;
 wire \soc/cpu/_03278_ ;
 wire \soc/cpu/_03279_ ;
 wire \soc/cpu/_03280_ ;
 wire \soc/cpu/_03281_ ;
 wire \soc/cpu/_03282_ ;
 wire \soc/cpu/_03283_ ;
 wire \soc/cpu/_03284_ ;
 wire \soc/cpu/_03285_ ;
 wire \soc/cpu/_03286_ ;
 wire \soc/cpu/_03287_ ;
 wire \soc/cpu/_03288_ ;
 wire \soc/cpu/_03289_ ;
 wire \soc/cpu/_03290_ ;
 wire \soc/cpu/_03291_ ;
 wire \soc/cpu/_03292_ ;
 wire \soc/cpu/_03293_ ;
 wire \soc/cpu/_03294_ ;
 wire \soc/cpu/_03295_ ;
 wire \soc/cpu/_03296_ ;
 wire \soc/cpu/_03297_ ;
 wire \soc/cpu/_03298_ ;
 wire \soc/cpu/_03299_ ;
 wire \soc/cpu/_03300_ ;
 wire net813;
 wire \soc/cpu/_03302_ ;
 wire \soc/cpu/_03303_ ;
 wire \soc/cpu/_03304_ ;
 wire \soc/cpu/_03305_ ;
 wire \soc/cpu/_03306_ ;
 wire \soc/cpu/_03307_ ;
 wire \soc/cpu/_03308_ ;
 wire \soc/cpu/_03309_ ;
 wire \soc/cpu/_03310_ ;
 wire \soc/cpu/_03311_ ;
 wire \soc/cpu/_03312_ ;
 wire \soc/cpu/_03313_ ;
 wire \soc/cpu/_03314_ ;
 wire \soc/cpu/_03315_ ;
 wire \soc/cpu/_03316_ ;
 wire \soc/cpu/_03317_ ;
 wire \soc/cpu/_03318_ ;
 wire \soc/cpu/_03319_ ;
 wire \soc/cpu/_03320_ ;
 wire \soc/cpu/_03321_ ;
 wire \soc/cpu/_03322_ ;
 wire \soc/cpu/_03323_ ;
 wire \soc/cpu/_03324_ ;
 wire \soc/cpu/_03325_ ;
 wire \soc/cpu/_03326_ ;
 wire \soc/cpu/_03327_ ;
 wire \soc/cpu/_03328_ ;
 wire net812;
 wire \soc/cpu/_03330_ ;
 wire \soc/cpu/_03331_ ;
 wire \soc/cpu/_03332_ ;
 wire \soc/cpu/_03333_ ;
 wire \soc/cpu/_03334_ ;
 wire \soc/cpu/_03335_ ;
 wire \soc/cpu/_03336_ ;
 wire \soc/cpu/_03337_ ;
 wire net811;
 wire net810;
 wire \soc/cpu/_03340_ ;
 wire \soc/cpu/_03341_ ;
 wire \soc/cpu/_03342_ ;
 wire \soc/cpu/_03343_ ;
 wire \soc/cpu/_03344_ ;
 wire net809;
 wire \soc/cpu/_03346_ ;
 wire \soc/cpu/_03347_ ;
 wire \soc/cpu/_03348_ ;
 wire \soc/cpu/_03349_ ;
 wire \soc/cpu/_03350_ ;
 wire \soc/cpu/_03351_ ;
 wire \soc/cpu/_03352_ ;
 wire \soc/cpu/_03353_ ;
 wire \soc/cpu/_03354_ ;
 wire \soc/cpu/_03355_ ;
 wire \soc/cpu/_03356_ ;
 wire \soc/cpu/_03357_ ;
 wire \soc/cpu/_03358_ ;
 wire \soc/cpu/_03359_ ;
 wire \soc/cpu/_03360_ ;
 wire net808;
 wire \soc/cpu/_03362_ ;
 wire \soc/cpu/_03363_ ;
 wire \soc/cpu/_03364_ ;
 wire \soc/cpu/_03365_ ;
 wire \soc/cpu/_03366_ ;
 wire \soc/cpu/_03367_ ;
 wire \soc/cpu/_03368_ ;
 wire \soc/cpu/_03369_ ;
 wire \soc/cpu/_03370_ ;
 wire \soc/cpu/_03371_ ;
 wire \soc/cpu/_03372_ ;
 wire \soc/cpu/_03373_ ;
 wire net807;
 wire net806;
 wire \soc/cpu/_03376_ ;
 wire \soc/cpu/_03377_ ;
 wire \soc/cpu/_03378_ ;
 wire \soc/cpu/_03379_ ;
 wire \soc/cpu/_03380_ ;
 wire \soc/cpu/_03381_ ;
 wire \soc/cpu/_03382_ ;
 wire \soc/cpu/_03383_ ;
 wire \soc/cpu/_03384_ ;
 wire \soc/cpu/_03385_ ;
 wire \soc/cpu/_03386_ ;
 wire \soc/cpu/_03387_ ;
 wire \soc/cpu/_03388_ ;
 wire \soc/cpu/_03389_ ;
 wire \soc/cpu/_03390_ ;
 wire \soc/cpu/_03391_ ;
 wire \soc/cpu/_03392_ ;
 wire \soc/cpu/_03393_ ;
 wire net805;
 wire \soc/cpu/_03395_ ;
 wire \soc/cpu/_03396_ ;
 wire \soc/cpu/_03397_ ;
 wire \soc/cpu/_03398_ ;
 wire \soc/cpu/_03399_ ;
 wire net804;
 wire net803;
 wire \soc/cpu/_03402_ ;
 wire \soc/cpu/_03403_ ;
 wire \soc/cpu/_03404_ ;
 wire \soc/cpu/_03405_ ;
 wire net802;
 wire \soc/cpu/_03407_ ;
 wire \soc/cpu/_03408_ ;
 wire \soc/cpu/_03409_ ;
 wire net801;
 wire \soc/cpu/_03411_ ;
 wire \soc/cpu/_03412_ ;
 wire net800;
 wire \soc/cpu/_03414_ ;
 wire net799;
 wire \soc/cpu/_03416_ ;
 wire \soc/cpu/_03417_ ;
 wire net798;
 wire \soc/cpu/_03419_ ;
 wire \soc/cpu/_03420_ ;
 wire net797;
 wire \soc/cpu/_03422_ ;
 wire \soc/cpu/_03423_ ;
 wire \soc/cpu/_03424_ ;
 wire \soc/cpu/_03425_ ;
 wire \soc/cpu/_03426_ ;
 wire \soc/cpu/_03427_ ;
 wire \soc/cpu/_03428_ ;
 wire \soc/cpu/_03429_ ;
 wire \soc/cpu/_03430_ ;
 wire \soc/cpu/_03431_ ;
 wire net796;
 wire net795;
 wire \soc/cpu/_03434_ ;
 wire \soc/cpu/_03435_ ;
 wire \soc/cpu/_03436_ ;
 wire \soc/cpu/_03437_ ;
 wire \soc/cpu/_03438_ ;
 wire \soc/cpu/_03439_ ;
 wire \soc/cpu/_03440_ ;
 wire \soc/cpu/_03441_ ;
 wire \soc/cpu/_03442_ ;
 wire \soc/cpu/_03443_ ;
 wire \soc/cpu/_03444_ ;
 wire net794;
 wire \soc/cpu/_03446_ ;
 wire net793;
 wire \soc/cpu/_03448_ ;
 wire \soc/cpu/_03449_ ;
 wire \soc/cpu/_03450_ ;
 wire \soc/cpu/_03451_ ;
 wire \soc/cpu/_03452_ ;
 wire \soc/cpu/_03453_ ;
 wire \soc/cpu/_03454_ ;
 wire \soc/cpu/_03455_ ;
 wire \soc/cpu/_03456_ ;
 wire \soc/cpu/_03457_ ;
 wire \soc/cpu/_03458_ ;
 wire \soc/cpu/_03459_ ;
 wire \soc/cpu/_03460_ ;
 wire \soc/cpu/_03461_ ;
 wire \soc/cpu/_03462_ ;
 wire \soc/cpu/_03463_ ;
 wire \soc/cpu/_03464_ ;
 wire \soc/cpu/_03465_ ;
 wire \soc/cpu/_03466_ ;
 wire \soc/cpu/_03467_ ;
 wire \soc/cpu/_03468_ ;
 wire \soc/cpu/_03469_ ;
 wire \soc/cpu/_03470_ ;
 wire \soc/cpu/_03471_ ;
 wire \soc/cpu/_03472_ ;
 wire \soc/cpu/_03473_ ;
 wire \soc/cpu/_03474_ ;
 wire \soc/cpu/_03475_ ;
 wire \soc/cpu/_03476_ ;
 wire net792;
 wire \soc/cpu/_03478_ ;
 wire \soc/cpu/_03479_ ;
 wire \soc/cpu/_03480_ ;
 wire \soc/cpu/_03481_ ;
 wire \soc/cpu/_03482_ ;
 wire \soc/cpu/_03483_ ;
 wire \soc/cpu/_03484_ ;
 wire \soc/cpu/_03485_ ;
 wire \soc/cpu/_03486_ ;
 wire \soc/cpu/_03487_ ;
 wire \soc/cpu/_03488_ ;
 wire \soc/cpu/_03489_ ;
 wire \soc/cpu/_03490_ ;
 wire \soc/cpu/_03491_ ;
 wire \soc/cpu/_03492_ ;
 wire net791;
 wire net790;
 wire net789;
 wire \soc/cpu/_03496_ ;
 wire \soc/cpu/_03497_ ;
 wire net788;
 wire net787;
 wire \soc/cpu/_03500_ ;
 wire net786;
 wire \soc/cpu/_03502_ ;
 wire \soc/cpu/_03503_ ;
 wire \soc/cpu/_03504_ ;
 wire \soc/cpu/_03505_ ;
 wire \soc/cpu/_03506_ ;
 wire \soc/cpu/_03507_ ;
 wire \soc/cpu/_03508_ ;
 wire \soc/cpu/_03509_ ;
 wire \soc/cpu/_03510_ ;
 wire \soc/cpu/_03511_ ;
 wire \soc/cpu/_03512_ ;
 wire \soc/cpu/_03513_ ;
 wire \soc/cpu/_03514_ ;
 wire \soc/cpu/_03515_ ;
 wire net785;
 wire net784;
 wire \soc/cpu/_03518_ ;
 wire net783;
 wire net782;
 wire \soc/cpu/_03521_ ;
 wire net781;
 wire net780;
 wire net779;
 wire net778;
 wire net777;
 wire \soc/cpu/_03527_ ;
 wire \soc/cpu/_03528_ ;
 wire \soc/cpu/_03529_ ;
 wire \soc/cpu/_03530_ ;
 wire \soc/cpu/_03531_ ;
 wire \soc/cpu/_03532_ ;
 wire \soc/cpu/_03533_ ;
 wire net776;
 wire \soc/cpu/_03535_ ;
 wire \soc/cpu/_03536_ ;
 wire \soc/cpu/_03537_ ;
 wire \soc/cpu/_03538_ ;
 wire \soc/cpu/_03539_ ;
 wire \soc/cpu/_03540_ ;
 wire \soc/cpu/_03541_ ;
 wire \soc/cpu/_03542_ ;
 wire \soc/cpu/_03543_ ;
 wire \soc/cpu/_03544_ ;
 wire \soc/cpu/_03545_ ;
 wire \soc/cpu/_03546_ ;
 wire \soc/cpu/_03547_ ;
 wire \soc/cpu/_03548_ ;
 wire \soc/cpu/_03549_ ;
 wire \soc/cpu/_03550_ ;
 wire \soc/cpu/_03551_ ;
 wire \soc/cpu/_03552_ ;
 wire \soc/cpu/_03553_ ;
 wire \soc/cpu/_03554_ ;
 wire \soc/cpu/_03555_ ;
 wire \soc/cpu/_03556_ ;
 wire \soc/cpu/_03557_ ;
 wire \soc/cpu/_03558_ ;
 wire \soc/cpu/_03559_ ;
 wire \soc/cpu/_03560_ ;
 wire \soc/cpu/_03561_ ;
 wire \soc/cpu/_03562_ ;
 wire \soc/cpu/_03563_ ;
 wire \soc/cpu/_03564_ ;
 wire \soc/cpu/_03565_ ;
 wire \soc/cpu/_03566_ ;
 wire \soc/cpu/_03567_ ;
 wire \soc/cpu/_03568_ ;
 wire \soc/cpu/_03569_ ;
 wire \soc/cpu/_03570_ ;
 wire \soc/cpu/_03571_ ;
 wire \soc/cpu/_03572_ ;
 wire \soc/cpu/_03573_ ;
 wire \soc/cpu/_03574_ ;
 wire \soc/cpu/_03575_ ;
 wire net775;
 wire \soc/cpu/_03577_ ;
 wire \soc/cpu/_03578_ ;
 wire \soc/cpu/_03579_ ;
 wire \soc/cpu/_03580_ ;
 wire \soc/cpu/_03581_ ;
 wire \soc/cpu/_03582_ ;
 wire \soc/cpu/_03583_ ;
 wire \soc/cpu/_03584_ ;
 wire \soc/cpu/_03585_ ;
 wire \soc/cpu/_03586_ ;
 wire \soc/cpu/_03587_ ;
 wire \soc/cpu/_03588_ ;
 wire \soc/cpu/_03589_ ;
 wire \soc/cpu/_03590_ ;
 wire \soc/cpu/_03591_ ;
 wire \soc/cpu/_03592_ ;
 wire \soc/cpu/_03593_ ;
 wire \soc/cpu/_03594_ ;
 wire \soc/cpu/_03595_ ;
 wire \soc/cpu/_03596_ ;
 wire \soc/cpu/_03597_ ;
 wire \soc/cpu/_03598_ ;
 wire \soc/cpu/_03599_ ;
 wire \soc/cpu/_03600_ ;
 wire \soc/cpu/_03601_ ;
 wire \soc/cpu/_03602_ ;
 wire \soc/cpu/_03603_ ;
 wire \soc/cpu/_03604_ ;
 wire \soc/cpu/_03605_ ;
 wire \soc/cpu/_03606_ ;
 wire \soc/cpu/_03607_ ;
 wire \soc/cpu/_03608_ ;
 wire \soc/cpu/_03609_ ;
 wire \soc/cpu/_03610_ ;
 wire \soc/cpu/_03611_ ;
 wire \soc/cpu/_03612_ ;
 wire \soc/cpu/_03613_ ;
 wire net774;
 wire \soc/cpu/_03615_ ;
 wire \soc/cpu/_03616_ ;
 wire \soc/cpu/_03617_ ;
 wire \soc/cpu/_03618_ ;
 wire \soc/cpu/_03619_ ;
 wire \soc/cpu/_03620_ ;
 wire \soc/cpu/_03621_ ;
 wire \soc/cpu/_03622_ ;
 wire \soc/cpu/_03623_ ;
 wire \soc/cpu/_03624_ ;
 wire \soc/cpu/_03625_ ;
 wire \soc/cpu/_03626_ ;
 wire \soc/cpu/_03627_ ;
 wire \soc/cpu/_03628_ ;
 wire \soc/cpu/_03629_ ;
 wire \soc/cpu/_03630_ ;
 wire \soc/cpu/_03631_ ;
 wire \soc/cpu/_03632_ ;
 wire \soc/cpu/_03633_ ;
 wire \soc/cpu/_03634_ ;
 wire \soc/cpu/_03635_ ;
 wire \soc/cpu/_03636_ ;
 wire \soc/cpu/_03637_ ;
 wire \soc/cpu/_03638_ ;
 wire \soc/cpu/_03639_ ;
 wire \soc/cpu/_03640_ ;
 wire \soc/cpu/_03641_ ;
 wire \soc/cpu/_03642_ ;
 wire \soc/cpu/_03643_ ;
 wire \soc/cpu/_03644_ ;
 wire \soc/cpu/_03645_ ;
 wire \soc/cpu/_03646_ ;
 wire \soc/cpu/_03647_ ;
 wire \soc/cpu/_03648_ ;
 wire \soc/cpu/_03649_ ;
 wire \soc/cpu/_03650_ ;
 wire \soc/cpu/_03651_ ;
 wire \soc/cpu/_03652_ ;
 wire \soc/cpu/_03653_ ;
 wire \soc/cpu/_03654_ ;
 wire \soc/cpu/_03655_ ;
 wire \soc/cpu/_03656_ ;
 wire \soc/cpu/_03657_ ;
 wire \soc/cpu/_03658_ ;
 wire \soc/cpu/_03659_ ;
 wire \soc/cpu/_03660_ ;
 wire \soc/cpu/_03661_ ;
 wire \soc/cpu/_03662_ ;
 wire \soc/cpu/_03663_ ;
 wire \soc/cpu/_03664_ ;
 wire \soc/cpu/_03665_ ;
 wire \soc/cpu/_03666_ ;
 wire \soc/cpu/_03667_ ;
 wire \soc/cpu/_03668_ ;
 wire \soc/cpu/_03669_ ;
 wire \soc/cpu/_03670_ ;
 wire \soc/cpu/_03671_ ;
 wire \soc/cpu/_03672_ ;
 wire \soc/cpu/_03673_ ;
 wire \soc/cpu/_03674_ ;
 wire \soc/cpu/_03675_ ;
 wire \soc/cpu/_03676_ ;
 wire \soc/cpu/_03677_ ;
 wire \soc/cpu/_03678_ ;
 wire \soc/cpu/_03679_ ;
 wire \soc/cpu/_03680_ ;
 wire \soc/cpu/_03681_ ;
 wire \soc/cpu/_03682_ ;
 wire net773;
 wire \soc/cpu/_03684_ ;
 wire \soc/cpu/_03685_ ;
 wire \soc/cpu/_03686_ ;
 wire \soc/cpu/_03687_ ;
 wire \soc/cpu/_03688_ ;
 wire \soc/cpu/_03689_ ;
 wire \soc/cpu/_03690_ ;
 wire \soc/cpu/_03691_ ;
 wire \soc/cpu/_03692_ ;
 wire \soc/cpu/_03693_ ;
 wire \soc/cpu/_03694_ ;
 wire \soc/cpu/_03695_ ;
 wire \soc/cpu/_03696_ ;
 wire \soc/cpu/_03697_ ;
 wire \soc/cpu/_03698_ ;
 wire \soc/cpu/_03699_ ;
 wire \soc/cpu/_03700_ ;
 wire \soc/cpu/_03701_ ;
 wire \soc/cpu/_03702_ ;
 wire \soc/cpu/_03703_ ;
 wire \soc/cpu/_03704_ ;
 wire \soc/cpu/_03705_ ;
 wire net772;
 wire net771;
 wire \soc/cpu/_03708_ ;
 wire \soc/cpu/_03709_ ;
 wire \soc/cpu/_03710_ ;
 wire \soc/cpu/_03711_ ;
 wire \soc/cpu/_03712_ ;
 wire \soc/cpu/_03713_ ;
 wire \soc/cpu/_03714_ ;
 wire \soc/cpu/_03715_ ;
 wire \soc/cpu/_03716_ ;
 wire \soc/cpu/_03717_ ;
 wire \soc/cpu/_03718_ ;
 wire \soc/cpu/_03719_ ;
 wire \soc/cpu/_03720_ ;
 wire \soc/cpu/_03721_ ;
 wire \soc/cpu/_03722_ ;
 wire \soc/cpu/_03723_ ;
 wire \soc/cpu/_03724_ ;
 wire \soc/cpu/_03725_ ;
 wire \soc/cpu/_03726_ ;
 wire \soc/cpu/_03727_ ;
 wire \soc/cpu/_03728_ ;
 wire \soc/cpu/_03729_ ;
 wire \soc/cpu/_03730_ ;
 wire \soc/cpu/_03731_ ;
 wire \soc/cpu/_03732_ ;
 wire \soc/cpu/_03733_ ;
 wire \soc/cpu/_03734_ ;
 wire \soc/cpu/_03735_ ;
 wire \soc/cpu/_03736_ ;
 wire \soc/cpu/_03737_ ;
 wire \soc/cpu/_03738_ ;
 wire \soc/cpu/_03739_ ;
 wire \soc/cpu/_03740_ ;
 wire \soc/cpu/_03741_ ;
 wire \soc/cpu/_03742_ ;
 wire \soc/cpu/_03743_ ;
 wire \soc/cpu/_03744_ ;
 wire \soc/cpu/_03745_ ;
 wire \soc/cpu/_03746_ ;
 wire \soc/cpu/_03747_ ;
 wire \soc/cpu/_03748_ ;
 wire \soc/cpu/_03749_ ;
 wire \soc/cpu/_03750_ ;
 wire \soc/cpu/_03751_ ;
 wire \soc/cpu/_03752_ ;
 wire \soc/cpu/_03753_ ;
 wire \soc/cpu/_03754_ ;
 wire \soc/cpu/_03755_ ;
 wire \soc/cpu/_03756_ ;
 wire \soc/cpu/_03757_ ;
 wire \soc/cpu/_03758_ ;
 wire \soc/cpu/_03759_ ;
 wire \soc/cpu/_03760_ ;
 wire \soc/cpu/_03761_ ;
 wire \soc/cpu/_03762_ ;
 wire \soc/cpu/_03763_ ;
 wire \soc/cpu/_03764_ ;
 wire \soc/cpu/_03765_ ;
 wire \soc/cpu/_03766_ ;
 wire \soc/cpu/_03767_ ;
 wire \soc/cpu/_03768_ ;
 wire \soc/cpu/_03769_ ;
 wire \soc/cpu/_03770_ ;
 wire \soc/cpu/_03771_ ;
 wire \soc/cpu/_03772_ ;
 wire \soc/cpu/_03773_ ;
 wire \soc/cpu/_03774_ ;
 wire \soc/cpu/_03775_ ;
 wire \soc/cpu/_03776_ ;
 wire \soc/cpu/_03777_ ;
 wire \soc/cpu/_03778_ ;
 wire \soc/cpu/_03779_ ;
 wire \soc/cpu/_03780_ ;
 wire \soc/cpu/_03781_ ;
 wire \soc/cpu/_03782_ ;
 wire \soc/cpu/_03783_ ;
 wire \soc/cpu/_03784_ ;
 wire \soc/cpu/_03785_ ;
 wire \soc/cpu/_03786_ ;
 wire \soc/cpu/_03787_ ;
 wire \soc/cpu/_03788_ ;
 wire \soc/cpu/_03789_ ;
 wire \soc/cpu/_03790_ ;
 wire \soc/cpu/_03791_ ;
 wire \soc/cpu/_03792_ ;
 wire \soc/cpu/_03793_ ;
 wire \soc/cpu/_03794_ ;
 wire \soc/cpu/_03795_ ;
 wire \soc/cpu/_03796_ ;
 wire \soc/cpu/_03797_ ;
 wire \soc/cpu/_03798_ ;
 wire \soc/cpu/_03799_ ;
 wire \soc/cpu/_03800_ ;
 wire \soc/cpu/_03801_ ;
 wire \soc/cpu/_03802_ ;
 wire \soc/cpu/_03803_ ;
 wire \soc/cpu/_03804_ ;
 wire \soc/cpu/_03805_ ;
 wire \soc/cpu/_03806_ ;
 wire \soc/cpu/_03807_ ;
 wire \soc/cpu/_03808_ ;
 wire \soc/cpu/_03809_ ;
 wire \soc/cpu/_03810_ ;
 wire \soc/cpu/_03811_ ;
 wire \soc/cpu/_03812_ ;
 wire \soc/cpu/_03813_ ;
 wire \soc/cpu/_03814_ ;
 wire \soc/cpu/_03815_ ;
 wire \soc/cpu/_03816_ ;
 wire \soc/cpu/_03817_ ;
 wire \soc/cpu/_03818_ ;
 wire \soc/cpu/_03819_ ;
 wire \soc/cpu/_03820_ ;
 wire \soc/cpu/_03821_ ;
 wire \soc/cpu/_03822_ ;
 wire \soc/cpu/_03823_ ;
 wire \soc/cpu/_03824_ ;
 wire \soc/cpu/_03825_ ;
 wire \soc/cpu/_03826_ ;
 wire \soc/cpu/_03827_ ;
 wire \soc/cpu/_03828_ ;
 wire \soc/cpu/_03829_ ;
 wire \soc/cpu/_03830_ ;
 wire \soc/cpu/_03831_ ;
 wire \soc/cpu/_03832_ ;
 wire \soc/cpu/_03833_ ;
 wire \soc/cpu/_03834_ ;
 wire \soc/cpu/_03835_ ;
 wire \soc/cpu/_03836_ ;
 wire \soc/cpu/_03837_ ;
 wire \soc/cpu/_03838_ ;
 wire \soc/cpu/_03839_ ;
 wire \soc/cpu/_03840_ ;
 wire \soc/cpu/_03841_ ;
 wire \soc/cpu/_03842_ ;
 wire \soc/cpu/_03843_ ;
 wire \soc/cpu/_03844_ ;
 wire \soc/cpu/_03845_ ;
 wire \soc/cpu/_03846_ ;
 wire \soc/cpu/_03847_ ;
 wire \soc/cpu/_03848_ ;
 wire \soc/cpu/_03849_ ;
 wire \soc/cpu/_03850_ ;
 wire \soc/cpu/_03851_ ;
 wire \soc/cpu/_03852_ ;
 wire \soc/cpu/_03853_ ;
 wire \soc/cpu/_03854_ ;
 wire \soc/cpu/_03855_ ;
 wire \soc/cpu/_03856_ ;
 wire \soc/cpu/_03857_ ;
 wire \soc/cpu/_03858_ ;
 wire \soc/cpu/_03859_ ;
 wire \soc/cpu/_03860_ ;
 wire \soc/cpu/_03861_ ;
 wire \soc/cpu/_03862_ ;
 wire \soc/cpu/_03863_ ;
 wire \soc/cpu/_03864_ ;
 wire \soc/cpu/_03865_ ;
 wire \soc/cpu/_03866_ ;
 wire \soc/cpu/_03867_ ;
 wire \soc/cpu/_03868_ ;
 wire \soc/cpu/_03869_ ;
 wire \soc/cpu/_03870_ ;
 wire \soc/cpu/_03871_ ;
 wire \soc/cpu/_03872_ ;
 wire \soc/cpu/_03873_ ;
 wire \soc/cpu/_03874_ ;
 wire \soc/cpu/_03875_ ;
 wire \soc/cpu/_03876_ ;
 wire \soc/cpu/_03877_ ;
 wire \soc/cpu/_03878_ ;
 wire \soc/cpu/_03879_ ;
 wire \soc/cpu/_03880_ ;
 wire \soc/cpu/_03881_ ;
 wire \soc/cpu/_03882_ ;
 wire \soc/cpu/_03883_ ;
 wire \soc/cpu/_03884_ ;
 wire \soc/cpu/_03885_ ;
 wire \soc/cpu/_03886_ ;
 wire \soc/cpu/_03887_ ;
 wire \soc/cpu/_03888_ ;
 wire \soc/cpu/_03889_ ;
 wire \soc/cpu/_03890_ ;
 wire \soc/cpu/_03891_ ;
 wire \soc/cpu/_03892_ ;
 wire \soc/cpu/_03893_ ;
 wire \soc/cpu/_03894_ ;
 wire \soc/cpu/_03895_ ;
 wire \soc/cpu/_03896_ ;
 wire \soc/cpu/_03897_ ;
 wire \soc/cpu/_03898_ ;
 wire \soc/cpu/_03899_ ;
 wire net770;
 wire \soc/cpu/_03901_ ;
 wire \soc/cpu/_03902_ ;
 wire \soc/cpu/_03903_ ;
 wire \soc/cpu/_03904_ ;
 wire \soc/cpu/_03905_ ;
 wire \soc/cpu/_03906_ ;
 wire \soc/cpu/_03907_ ;
 wire \soc/cpu/_03908_ ;
 wire \soc/cpu/_03909_ ;
 wire \soc/cpu/_03910_ ;
 wire \soc/cpu/_03911_ ;
 wire \soc/cpu/_03912_ ;
 wire \soc/cpu/_03913_ ;
 wire \soc/cpu/_03914_ ;
 wire \soc/cpu/_03915_ ;
 wire \soc/cpu/_03916_ ;
 wire \soc/cpu/_03917_ ;
 wire \soc/cpu/_03918_ ;
 wire \soc/cpu/_03919_ ;
 wire \soc/cpu/_03920_ ;
 wire \soc/cpu/_03921_ ;
 wire \soc/cpu/_03922_ ;
 wire \soc/cpu/_03923_ ;
 wire \soc/cpu/_03924_ ;
 wire \soc/cpu/_03925_ ;
 wire \soc/cpu/_03926_ ;
 wire \soc/cpu/_03927_ ;
 wire \soc/cpu/_03928_ ;
 wire \soc/cpu/_03929_ ;
 wire \soc/cpu/_03930_ ;
 wire \soc/cpu/_03931_ ;
 wire \soc/cpu/_03932_ ;
 wire \soc/cpu/_03933_ ;
 wire \soc/cpu/_03934_ ;
 wire \soc/cpu/_03935_ ;
 wire \soc/cpu/_03936_ ;
 wire \soc/cpu/_03937_ ;
 wire \soc/cpu/_03938_ ;
 wire \soc/cpu/_03939_ ;
 wire \soc/cpu/_03940_ ;
 wire \soc/cpu/_03941_ ;
 wire \soc/cpu/_03942_ ;
 wire \soc/cpu/_03943_ ;
 wire \soc/cpu/_03944_ ;
 wire \soc/cpu/_03945_ ;
 wire \soc/cpu/_03946_ ;
 wire net769;
 wire net768;
 wire \soc/cpu/_03949_ ;
 wire net767;
 wire \soc/cpu/_03951_ ;
 wire \soc/cpu/_03952_ ;
 wire \soc/cpu/_03953_ ;
 wire \soc/cpu/_03954_ ;
 wire \soc/cpu/_03955_ ;
 wire \soc/cpu/_03956_ ;
 wire \soc/cpu/_03957_ ;
 wire net766;
 wire \soc/cpu/_03959_ ;
 wire \soc/cpu/_03960_ ;
 wire net765;
 wire \soc/cpu/_03962_ ;
 wire net764;
 wire \soc/cpu/_03964_ ;
 wire \soc/cpu/_03965_ ;
 wire \soc/cpu/_03966_ ;
 wire \soc/cpu/_03967_ ;
 wire \soc/cpu/_03968_ ;
 wire \soc/cpu/_03969_ ;
 wire \soc/cpu/_03970_ ;
 wire net763;
 wire \soc/cpu/_03972_ ;
 wire \soc/cpu/_03973_ ;
 wire net762;
 wire \soc/cpu/_03975_ ;
 wire net761;
 wire \soc/cpu/_03977_ ;
 wire \soc/cpu/_03978_ ;
 wire \soc/cpu/_03979_ ;
 wire \soc/cpu/_03980_ ;
 wire \soc/cpu/_03981_ ;
 wire \soc/cpu/_03982_ ;
 wire \soc/cpu/_03983_ ;
 wire \soc/cpu/_03984_ ;
 wire \soc/cpu/_03985_ ;
 wire \soc/cpu/_03986_ ;
 wire net760;
 wire \soc/cpu/_03988_ ;
 wire \soc/cpu/_03989_ ;
 wire \soc/cpu/_03990_ ;
 wire \soc/cpu/_03991_ ;
 wire \soc/cpu/_03992_ ;
 wire \soc/cpu/_03993_ ;
 wire \soc/cpu/_03994_ ;
 wire \soc/cpu/_03995_ ;
 wire \soc/cpu/_03996_ ;
 wire \soc/cpu/_03997_ ;
 wire \soc/cpu/_03998_ ;
 wire \soc/cpu/_03999_ ;
 wire \soc/cpu/_04000_ ;
 wire \soc/cpu/_04001_ ;
 wire \soc/cpu/_04002_ ;
 wire \soc/cpu/_04003_ ;
 wire \soc/cpu/_04004_ ;
 wire \soc/cpu/_04005_ ;
 wire \soc/cpu/_04006_ ;
 wire \soc/cpu/_04007_ ;
 wire \soc/cpu/_04008_ ;
 wire \soc/cpu/_04009_ ;
 wire \soc/cpu/_04010_ ;
 wire \soc/cpu/_04011_ ;
 wire \soc/cpu/_04012_ ;
 wire \soc/cpu/_04013_ ;
 wire \soc/cpu/_04014_ ;
 wire \soc/cpu/_04015_ ;
 wire \soc/cpu/_04016_ ;
 wire \soc/cpu/_04017_ ;
 wire \soc/cpu/_04018_ ;
 wire \soc/cpu/_04019_ ;
 wire \soc/cpu/_04020_ ;
 wire \soc/cpu/_04021_ ;
 wire \soc/cpu/_04022_ ;
 wire \soc/cpu/_04023_ ;
 wire \soc/cpu/_04024_ ;
 wire net759;
 wire \soc/cpu/_04026_ ;
 wire \soc/cpu/_04027_ ;
 wire \soc/cpu/_04028_ ;
 wire net758;
 wire \soc/cpu/_04030_ ;
 wire \soc/cpu/_04031_ ;
 wire \soc/cpu/_04032_ ;
 wire \soc/cpu/_04033_ ;
 wire \soc/cpu/_04034_ ;
 wire \soc/cpu/_04035_ ;
 wire \soc/cpu/_04036_ ;
 wire \soc/cpu/_04037_ ;
 wire \soc/cpu/_04038_ ;
 wire \soc/cpu/_04039_ ;
 wire \soc/cpu/_04040_ ;
 wire \soc/cpu/_04041_ ;
 wire \soc/cpu/_04042_ ;
 wire \soc/cpu/_04043_ ;
 wire \soc/cpu/_04044_ ;
 wire \soc/cpu/_04045_ ;
 wire \soc/cpu/_04046_ ;
 wire \soc/cpu/_04047_ ;
 wire \soc/cpu/_04048_ ;
 wire \soc/cpu/_04049_ ;
 wire \soc/cpu/_04050_ ;
 wire \soc/cpu/_04051_ ;
 wire \soc/cpu/_04052_ ;
 wire \soc/cpu/_04053_ ;
 wire \soc/cpu/_04054_ ;
 wire \soc/cpu/_04055_ ;
 wire \soc/cpu/_04056_ ;
 wire \soc/cpu/_04057_ ;
 wire \soc/cpu/_04058_ ;
 wire \soc/cpu/_04059_ ;
 wire \soc/cpu/_04060_ ;
 wire \soc/cpu/_04061_ ;
 wire net757;
 wire \soc/cpu/_04063_ ;
 wire \soc/cpu/_04064_ ;
 wire net756;
 wire \soc/cpu/_04066_ ;
 wire \soc/cpu/_04067_ ;
 wire \soc/cpu/_04068_ ;
 wire \soc/cpu/_04069_ ;
 wire \soc/cpu/_04070_ ;
 wire \soc/cpu/_04071_ ;
 wire \soc/cpu/_04072_ ;
 wire \soc/cpu/_04073_ ;
 wire \soc/cpu/_04074_ ;
 wire \soc/cpu/_04075_ ;
 wire \soc/cpu/_04076_ ;
 wire \soc/cpu/_04077_ ;
 wire \soc/cpu/_04078_ ;
 wire \soc/cpu/_04079_ ;
 wire \soc/cpu/_04080_ ;
 wire \soc/cpu/_04081_ ;
 wire \soc/cpu/_04082_ ;
 wire \soc/cpu/_04083_ ;
 wire \soc/cpu/_04084_ ;
 wire \soc/cpu/_04085_ ;
 wire \soc/cpu/_04086_ ;
 wire \soc/cpu/_04087_ ;
 wire \soc/cpu/_04088_ ;
 wire \soc/cpu/_04089_ ;
 wire \soc/cpu/_04090_ ;
 wire \soc/cpu/_04091_ ;
 wire \soc/cpu/_04092_ ;
 wire \soc/cpu/_04093_ ;
 wire \soc/cpu/_04094_ ;
 wire \soc/cpu/_04095_ ;
 wire \soc/cpu/_04096_ ;
 wire \soc/cpu/_04097_ ;
 wire \soc/cpu/_04098_ ;
 wire \soc/cpu/_04099_ ;
 wire \soc/cpu/_04100_ ;
 wire \soc/cpu/_04101_ ;
 wire \soc/cpu/_04102_ ;
 wire \soc/cpu/_04103_ ;
 wire \soc/cpu/_04104_ ;
 wire \soc/cpu/_04105_ ;
 wire \soc/cpu/_04106_ ;
 wire \soc/cpu/_04107_ ;
 wire \soc/cpu/_04108_ ;
 wire \soc/cpu/_04109_ ;
 wire net755;
 wire \soc/cpu/_04111_ ;
 wire \soc/cpu/_04112_ ;
 wire \soc/cpu/_04113_ ;
 wire \soc/cpu/_04114_ ;
 wire net754;
 wire \soc/cpu/_04116_ ;
 wire net753;
 wire \soc/cpu/_04118_ ;
 wire \soc/cpu/_04119_ ;
 wire \soc/cpu/_04120_ ;
 wire \soc/cpu/_04121_ ;
 wire \soc/cpu/_04122_ ;
 wire \soc/cpu/_04123_ ;
 wire \soc/cpu/_04124_ ;
 wire \soc/cpu/_04125_ ;
 wire \soc/cpu/_04126_ ;
 wire \soc/cpu/_04127_ ;
 wire \soc/cpu/_04128_ ;
 wire net752;
 wire \soc/cpu/_04130_ ;
 wire \soc/cpu/_04131_ ;
 wire net751;
 wire \soc/cpu/_04133_ ;
 wire \soc/cpu/_04134_ ;
 wire \soc/cpu/_04135_ ;
 wire \soc/cpu/_04136_ ;
 wire \soc/cpu/_04137_ ;
 wire \soc/cpu/_04138_ ;
 wire \soc/cpu/_04139_ ;
 wire \soc/cpu/_04140_ ;
 wire \soc/cpu/_04141_ ;
 wire net750;
 wire \soc/cpu/_04143_ ;
 wire \soc/cpu/_04144_ ;
 wire \soc/cpu/_04145_ ;
 wire \soc/cpu/_04146_ ;
 wire \soc/cpu/_04147_ ;
 wire \soc/cpu/_04148_ ;
 wire \soc/cpu/_04149_ ;
 wire \soc/cpu/_04150_ ;
 wire \soc/cpu/_04151_ ;
 wire \soc/cpu/_04152_ ;
 wire \soc/cpu/_04153_ ;
 wire \soc/cpu/_04154_ ;
 wire \soc/cpu/_04155_ ;
 wire \soc/cpu/_04156_ ;
 wire \soc/cpu/_04157_ ;
 wire net749;
 wire \soc/cpu/_04159_ ;
 wire \soc/cpu/_04160_ ;
 wire \soc/cpu/_04161_ ;
 wire \soc/cpu/_04162_ ;
 wire \soc/cpu/_04163_ ;
 wire \soc/cpu/_04164_ ;
 wire \soc/cpu/_04165_ ;
 wire \soc/cpu/_04166_ ;
 wire \soc/cpu/_04167_ ;
 wire \soc/cpu/_04168_ ;
 wire \soc/cpu/_04169_ ;
 wire \soc/cpu/_04170_ ;
 wire \soc/cpu/_04171_ ;
 wire \soc/cpu/_04172_ ;
 wire \soc/cpu/_04173_ ;
 wire \soc/cpu/_04174_ ;
 wire \soc/cpu/_04175_ ;
 wire \soc/cpu/_04176_ ;
 wire \soc/cpu/_04177_ ;
 wire \soc/cpu/_04178_ ;
 wire \soc/cpu/_04179_ ;
 wire \soc/cpu/_04180_ ;
 wire \soc/cpu/_04181_ ;
 wire \soc/cpu/_04182_ ;
 wire \soc/cpu/_04183_ ;
 wire \soc/cpu/_04184_ ;
 wire \soc/cpu/_04185_ ;
 wire \soc/cpu/_04186_ ;
 wire \soc/cpu/_04187_ ;
 wire \soc/cpu/_04188_ ;
 wire \soc/cpu/_04189_ ;
 wire \soc/cpu/_04190_ ;
 wire \soc/cpu/_04191_ ;
 wire \soc/cpu/_04192_ ;
 wire \soc/cpu/_04193_ ;
 wire \soc/cpu/_04194_ ;
 wire \soc/cpu/_04195_ ;
 wire \soc/cpu/_04196_ ;
 wire \soc/cpu/_04197_ ;
 wire \soc/cpu/_04198_ ;
 wire \soc/cpu/_04199_ ;
 wire \soc/cpu/_04200_ ;
 wire \soc/cpu/_04201_ ;
 wire \soc/cpu/_04202_ ;
 wire \soc/cpu/_04203_ ;
 wire net748;
 wire \soc/cpu/_04205_ ;
 wire \soc/cpu/_04206_ ;
 wire \soc/cpu/_04207_ ;
 wire \soc/cpu/_04208_ ;
 wire \soc/cpu/_04209_ ;
 wire \soc/cpu/_04210_ ;
 wire \soc/cpu/_04211_ ;
 wire \soc/cpu/_04212_ ;
 wire \soc/cpu/_04213_ ;
 wire \soc/cpu/_04214_ ;
 wire \soc/cpu/_04215_ ;
 wire \soc/cpu/_04216_ ;
 wire \soc/cpu/_04217_ ;
 wire \soc/cpu/_04218_ ;
 wire \soc/cpu/_04219_ ;
 wire \soc/cpu/_04220_ ;
 wire \soc/cpu/_04221_ ;
 wire \soc/cpu/_04222_ ;
 wire net747;
 wire net746;
 wire \soc/cpu/_04225_ ;
 wire \soc/cpu/_04226_ ;
 wire \soc/cpu/_04227_ ;
 wire \soc/cpu/_04228_ ;
 wire net745;
 wire \soc/cpu/_04230_ ;
 wire \soc/cpu/_04231_ ;
 wire \soc/cpu/_04232_ ;
 wire \soc/cpu/_04233_ ;
 wire \soc/cpu/_04234_ ;
 wire \soc/cpu/_04235_ ;
 wire \soc/cpu/_04236_ ;
 wire \soc/cpu/_04237_ ;
 wire \soc/cpu/_04238_ ;
 wire \soc/cpu/_04239_ ;
 wire \soc/cpu/_04240_ ;
 wire \soc/cpu/_04241_ ;
 wire \soc/cpu/_04242_ ;
 wire \soc/cpu/_04243_ ;
 wire \soc/cpu/_04244_ ;
 wire \soc/cpu/_04245_ ;
 wire \soc/cpu/_04246_ ;
 wire \soc/cpu/_04247_ ;
 wire \soc/cpu/_04248_ ;
 wire \soc/cpu/_04249_ ;
 wire \soc/cpu/_04250_ ;
 wire \soc/cpu/_04251_ ;
 wire net744;
 wire \soc/cpu/_04253_ ;
 wire \soc/cpu/_04254_ ;
 wire \soc/cpu/_04255_ ;
 wire \soc/cpu/_04256_ ;
 wire \soc/cpu/_04257_ ;
 wire \soc/cpu/_04258_ ;
 wire \soc/cpu/_04259_ ;
 wire \soc/cpu/_04260_ ;
 wire \soc/cpu/_04261_ ;
 wire \soc/cpu/_04262_ ;
 wire \soc/cpu/_04263_ ;
 wire \soc/cpu/_04264_ ;
 wire \soc/cpu/_04265_ ;
 wire \soc/cpu/_04266_ ;
 wire \soc/cpu/_04267_ ;
 wire \soc/cpu/_04268_ ;
 wire \soc/cpu/_04269_ ;
 wire \soc/cpu/_04270_ ;
 wire \soc/cpu/_04271_ ;
 wire \soc/cpu/_04272_ ;
 wire \soc/cpu/_04273_ ;
 wire \soc/cpu/_04274_ ;
 wire \soc/cpu/_04275_ ;
 wire \soc/cpu/_04276_ ;
 wire \soc/cpu/_04277_ ;
 wire \soc/cpu/_04278_ ;
 wire \soc/cpu/_04279_ ;
 wire \soc/cpu/_04280_ ;
 wire \soc/cpu/_04281_ ;
 wire \soc/cpu/_04282_ ;
 wire \soc/cpu/_04283_ ;
 wire \soc/cpu/_04284_ ;
 wire \soc/cpu/_04285_ ;
 wire \soc/cpu/_04286_ ;
 wire \soc/cpu/_04287_ ;
 wire \soc/cpu/_04288_ ;
 wire \soc/cpu/_04289_ ;
 wire \soc/cpu/_04290_ ;
 wire \soc/cpu/_04291_ ;
 wire \soc/cpu/_04292_ ;
 wire \soc/cpu/_04293_ ;
 wire net743;
 wire \soc/cpu/_04295_ ;
 wire \soc/cpu/_04296_ ;
 wire \soc/cpu/_04297_ ;
 wire \soc/cpu/_04298_ ;
 wire \soc/cpu/_04299_ ;
 wire \soc/cpu/_04300_ ;
 wire \soc/cpu/_04301_ ;
 wire \soc/cpu/_04302_ ;
 wire \soc/cpu/_04303_ ;
 wire \soc/cpu/_04304_ ;
 wire \soc/cpu/_04305_ ;
 wire \soc/cpu/_04306_ ;
 wire \soc/cpu/_04307_ ;
 wire \soc/cpu/_04308_ ;
 wire \soc/cpu/_04309_ ;
 wire \soc/cpu/_04310_ ;
 wire \soc/cpu/_04311_ ;
 wire \soc/cpu/_04312_ ;
 wire \soc/cpu/_04313_ ;
 wire \soc/cpu/_04314_ ;
 wire \soc/cpu/_04315_ ;
 wire \soc/cpu/_04316_ ;
 wire \soc/cpu/_04317_ ;
 wire \soc/cpu/_04318_ ;
 wire \soc/cpu/_04319_ ;
 wire \soc/cpu/_04320_ ;
 wire \soc/cpu/_04321_ ;
 wire \soc/cpu/_04322_ ;
 wire \soc/cpu/_04323_ ;
 wire \soc/cpu/_04324_ ;
 wire \soc/cpu/_04325_ ;
 wire \soc/cpu/_04326_ ;
 wire \soc/cpu/_04327_ ;
 wire \soc/cpu/_04328_ ;
 wire \soc/cpu/_04329_ ;
 wire net742;
 wire \soc/cpu/_04331_ ;
 wire \soc/cpu/_04332_ ;
 wire \soc/cpu/_04333_ ;
 wire \soc/cpu/_04334_ ;
 wire \soc/cpu/_04335_ ;
 wire \soc/cpu/_04336_ ;
 wire \soc/cpu/_04337_ ;
 wire \soc/cpu/_04338_ ;
 wire \soc/cpu/_04339_ ;
 wire \soc/cpu/_04340_ ;
 wire \soc/cpu/_04341_ ;
 wire \soc/cpu/_04342_ ;
 wire \soc/cpu/_04343_ ;
 wire \soc/cpu/_04344_ ;
 wire \soc/cpu/_04345_ ;
 wire \soc/cpu/_04346_ ;
 wire \soc/cpu/_04347_ ;
 wire \soc/cpu/_04348_ ;
 wire \soc/cpu/_04349_ ;
 wire \soc/cpu/_04350_ ;
 wire \soc/cpu/_04351_ ;
 wire \soc/cpu/_04352_ ;
 wire \soc/cpu/_04353_ ;
 wire \soc/cpu/_04354_ ;
 wire \soc/cpu/_04355_ ;
 wire \soc/cpu/_04356_ ;
 wire \soc/cpu/_04357_ ;
 wire \soc/cpu/_04358_ ;
 wire \soc/cpu/_04359_ ;
 wire \soc/cpu/_04360_ ;
 wire \soc/cpu/_04361_ ;
 wire \soc/cpu/_04362_ ;
 wire \soc/cpu/_04363_ ;
 wire \soc/cpu/_04364_ ;
 wire \soc/cpu/_04365_ ;
 wire \soc/cpu/_04366_ ;
 wire \soc/cpu/_04367_ ;
 wire \soc/cpu/_04368_ ;
 wire \soc/cpu/_04369_ ;
 wire \soc/cpu/_04370_ ;
 wire \soc/cpu/_04371_ ;
 wire \soc/cpu/_04372_ ;
 wire \soc/cpu/_04373_ ;
 wire \soc/cpu/_04374_ ;
 wire \soc/cpu/_04375_ ;
 wire \soc/cpu/_04376_ ;
 wire \soc/cpu/_04377_ ;
 wire \soc/cpu/_04378_ ;
 wire \soc/cpu/_04379_ ;
 wire \soc/cpu/_04380_ ;
 wire \soc/cpu/_04381_ ;
 wire \soc/cpu/_04382_ ;
 wire \soc/cpu/_04383_ ;
 wire \soc/cpu/_04384_ ;
 wire \soc/cpu/_04385_ ;
 wire \soc/cpu/_04386_ ;
 wire \soc/cpu/_04387_ ;
 wire \soc/cpu/_04388_ ;
 wire \soc/cpu/_04389_ ;
 wire \soc/cpu/_04390_ ;
 wire \soc/cpu/_04391_ ;
 wire \soc/cpu/_04392_ ;
 wire \soc/cpu/_04393_ ;
 wire \soc/cpu/_04394_ ;
 wire \soc/cpu/_04395_ ;
 wire \soc/cpu/_04396_ ;
 wire \soc/cpu/_04397_ ;
 wire \soc/cpu/_04398_ ;
 wire \soc/cpu/_04399_ ;
 wire \soc/cpu/_04400_ ;
 wire \soc/cpu/_04401_ ;
 wire \soc/cpu/_04402_ ;
 wire \soc/cpu/_04403_ ;
 wire \soc/cpu/_04404_ ;
 wire net741;
 wire \soc/cpu/_04406_ ;
 wire \soc/cpu/_04407_ ;
 wire \soc/cpu/_04408_ ;
 wire \soc/cpu/_04409_ ;
 wire \soc/cpu/_04410_ ;
 wire \soc/cpu/_04411_ ;
 wire \soc/cpu/_04412_ ;
 wire \soc/cpu/_04413_ ;
 wire \soc/cpu/_04414_ ;
 wire \soc/cpu/_04415_ ;
 wire \soc/cpu/_04416_ ;
 wire \soc/cpu/_04417_ ;
 wire \soc/cpu/_04418_ ;
 wire \soc/cpu/_04419_ ;
 wire \soc/cpu/_04420_ ;
 wire net740;
 wire \soc/cpu/_04422_ ;
 wire \soc/cpu/_04423_ ;
 wire \soc/cpu/_04424_ ;
 wire \soc/cpu/_04425_ ;
 wire \soc/cpu/_04426_ ;
 wire \soc/cpu/_04427_ ;
 wire \soc/cpu/_04428_ ;
 wire \soc/cpu/_04429_ ;
 wire \soc/cpu/_04430_ ;
 wire \soc/cpu/_04431_ ;
 wire \soc/cpu/_04432_ ;
 wire \soc/cpu/_04433_ ;
 wire \soc/cpu/_04434_ ;
 wire \soc/cpu/_04435_ ;
 wire \soc/cpu/_04436_ ;
 wire \soc/cpu/_04437_ ;
 wire \soc/cpu/_04438_ ;
 wire \soc/cpu/_04439_ ;
 wire \soc/cpu/_04440_ ;
 wire \soc/cpu/_04441_ ;
 wire \soc/cpu/_04442_ ;
 wire \soc/cpu/_04443_ ;
 wire \soc/cpu/_04444_ ;
 wire \soc/cpu/_04445_ ;
 wire \soc/cpu/_04446_ ;
 wire \soc/cpu/_04447_ ;
 wire \soc/cpu/_04448_ ;
 wire \soc/cpu/_04449_ ;
 wire \soc/cpu/_04450_ ;
 wire \soc/cpu/_04451_ ;
 wire \soc/cpu/_04452_ ;
 wire \soc/cpu/_04453_ ;
 wire \soc/cpu/_04454_ ;
 wire \soc/cpu/_04455_ ;
 wire \soc/cpu/_04456_ ;
 wire \soc/cpu/_04457_ ;
 wire \soc/cpu/_04458_ ;
 wire \soc/cpu/_04459_ ;
 wire \soc/cpu/_04460_ ;
 wire \soc/cpu/_04461_ ;
 wire \soc/cpu/_04462_ ;
 wire \soc/cpu/_04463_ ;
 wire \soc/cpu/_04464_ ;
 wire \soc/cpu/_04465_ ;
 wire \soc/cpu/_04466_ ;
 wire \soc/cpu/_04467_ ;
 wire \soc/cpu/_04468_ ;
 wire \soc/cpu/_04469_ ;
 wire \soc/cpu/_04470_ ;
 wire \soc/cpu/_04471_ ;
 wire \soc/cpu/_04472_ ;
 wire \soc/cpu/_04473_ ;
 wire \soc/cpu/_04474_ ;
 wire \soc/cpu/_04475_ ;
 wire \soc/cpu/_04476_ ;
 wire \soc/cpu/_04477_ ;
 wire \soc/cpu/_04478_ ;
 wire \soc/cpu/_04479_ ;
 wire \soc/cpu/_04480_ ;
 wire \soc/cpu/_04481_ ;
 wire \soc/cpu/_04482_ ;
 wire \soc/cpu/_04483_ ;
 wire \soc/cpu/_04484_ ;
 wire \soc/cpu/_04485_ ;
 wire \soc/cpu/_04486_ ;
 wire \soc/cpu/_04487_ ;
 wire \soc/cpu/_04488_ ;
 wire \soc/cpu/_04489_ ;
 wire \soc/cpu/_04490_ ;
 wire \soc/cpu/_04491_ ;
 wire \soc/cpu/_04492_ ;
 wire \soc/cpu/_04493_ ;
 wire \soc/cpu/_04494_ ;
 wire \soc/cpu/_04495_ ;
 wire \soc/cpu/_04496_ ;
 wire \soc/cpu/_04497_ ;
 wire \soc/cpu/_04498_ ;
 wire \soc/cpu/_04499_ ;
 wire \soc/cpu/_04500_ ;
 wire \soc/cpu/_04501_ ;
 wire \soc/cpu/_04502_ ;
 wire \soc/cpu/_04503_ ;
 wire \soc/cpu/_04504_ ;
 wire \soc/cpu/_04505_ ;
 wire \soc/cpu/_04506_ ;
 wire \soc/cpu/_04507_ ;
 wire \soc/cpu/_04508_ ;
 wire \soc/cpu/_04509_ ;
 wire \soc/cpu/_04510_ ;
 wire \soc/cpu/_04511_ ;
 wire \soc/cpu/_04512_ ;
 wire \soc/cpu/_04513_ ;
 wire \soc/cpu/_04514_ ;
 wire \soc/cpu/_04515_ ;
 wire \soc/cpu/_04516_ ;
 wire \soc/cpu/_04517_ ;
 wire \soc/cpu/_04518_ ;
 wire \soc/cpu/_04519_ ;
 wire \soc/cpu/_04520_ ;
 wire \soc/cpu/_04521_ ;
 wire \soc/cpu/_04522_ ;
 wire \soc/cpu/_04523_ ;
 wire \soc/cpu/_04524_ ;
 wire \soc/cpu/_04525_ ;
 wire \soc/cpu/_04526_ ;
 wire \soc/cpu/_04527_ ;
 wire \soc/cpu/_04528_ ;
 wire \soc/cpu/_04529_ ;
 wire \soc/cpu/_04530_ ;
 wire \soc/cpu/_04531_ ;
 wire \soc/cpu/_04532_ ;
 wire \soc/cpu/_04533_ ;
 wire \soc/cpu/_04534_ ;
 wire \soc/cpu/_04535_ ;
 wire \soc/cpu/_04536_ ;
 wire \soc/cpu/_04537_ ;
 wire \soc/cpu/_04538_ ;
 wire \soc/cpu/_04539_ ;
 wire \soc/cpu/_04540_ ;
 wire \soc/cpu/_04541_ ;
 wire \soc/cpu/_04542_ ;
 wire \soc/cpu/_04543_ ;
 wire \soc/cpu/_04544_ ;
 wire \soc/cpu/_04545_ ;
 wire \soc/cpu/_04546_ ;
 wire \soc/cpu/_04547_ ;
 wire \soc/cpu/_04548_ ;
 wire \soc/cpu/_04549_ ;
 wire \soc/cpu/_04550_ ;
 wire \soc/cpu/_04551_ ;
 wire \soc/cpu/_04552_ ;
 wire \soc/cpu/_04553_ ;
 wire \soc/cpu/_04554_ ;
 wire \soc/cpu/_04555_ ;
 wire \soc/cpu/_04556_ ;
 wire \soc/cpu/_04557_ ;
 wire \soc/cpu/_04558_ ;
 wire \soc/cpu/_04559_ ;
 wire \soc/cpu/_04560_ ;
 wire \soc/cpu/_04561_ ;
 wire \soc/cpu/_04562_ ;
 wire \soc/cpu/_04563_ ;
 wire \soc/cpu/_04564_ ;
 wire \soc/cpu/_04565_ ;
 wire \soc/cpu/_04566_ ;
 wire \soc/cpu/_04567_ ;
 wire \soc/cpu/_04568_ ;
 wire \soc/cpu/_04569_ ;
 wire \soc/cpu/_04570_ ;
 wire \soc/cpu/_04571_ ;
 wire net739;
 wire net738;
 wire \soc/cpu/_04574_ ;
 wire \soc/cpu/_04575_ ;
 wire \soc/cpu/_04576_ ;
 wire net737;
 wire net736;
 wire \soc/cpu/_04579_ ;
 wire net735;
 wire \soc/cpu/_04581_ ;
 wire \soc/cpu/_04582_ ;
 wire \soc/cpu/_04583_ ;
 wire \soc/cpu/_04584_ ;
 wire \soc/cpu/_04585_ ;
 wire \soc/cpu/_04586_ ;
 wire \soc/cpu/_04587_ ;
 wire net734;
 wire \soc/cpu/_04589_ ;
 wire \soc/cpu/_04590_ ;
 wire \soc/cpu/_04591_ ;
 wire \soc/cpu/_04592_ ;
 wire \soc/cpu/_04593_ ;
 wire \soc/cpu/_04594_ ;
 wire \soc/cpu/_04595_ ;
 wire \soc/cpu/_04596_ ;
 wire \soc/cpu/_04597_ ;
 wire \soc/cpu/_04598_ ;
 wire \soc/cpu/_04599_ ;
 wire \soc/cpu/_04600_ ;
 wire \soc/cpu/_04601_ ;
 wire \soc/cpu/_04602_ ;
 wire \soc/cpu/_04603_ ;
 wire \soc/cpu/_04604_ ;
 wire \soc/cpu/_04605_ ;
 wire \soc/cpu/_04606_ ;
 wire \soc/cpu/_04607_ ;
 wire \soc/cpu/_04608_ ;
 wire \soc/cpu/_04609_ ;
 wire \soc/cpu/_04610_ ;
 wire \soc/cpu/_04611_ ;
 wire \soc/cpu/_04612_ ;
 wire \soc/cpu/_04613_ ;
 wire \soc/cpu/_04614_ ;
 wire \soc/cpu/_04615_ ;
 wire \soc/cpu/_04616_ ;
 wire \soc/cpu/_04617_ ;
 wire \soc/cpu/_04618_ ;
 wire \soc/cpu/_04619_ ;
 wire \soc/cpu/_04620_ ;
 wire \soc/cpu/_04621_ ;
 wire \soc/cpu/_04622_ ;
 wire \soc/cpu/_04623_ ;
 wire \soc/cpu/_04624_ ;
 wire \soc/cpu/_04625_ ;
 wire \soc/cpu/_04626_ ;
 wire \soc/cpu/_04627_ ;
 wire net733;
 wire \soc/cpu/_04629_ ;
 wire \soc/cpu/_04630_ ;
 wire \soc/cpu/_04631_ ;
 wire \soc/cpu/_04632_ ;
 wire \soc/cpu/_04633_ ;
 wire \soc/cpu/_04634_ ;
 wire \soc/cpu/_04635_ ;
 wire \soc/cpu/_04636_ ;
 wire \soc/cpu/_04637_ ;
 wire \soc/cpu/_04638_ ;
 wire \soc/cpu/_04639_ ;
 wire \soc/cpu/_04640_ ;
 wire \soc/cpu/_04641_ ;
 wire \soc/cpu/_04642_ ;
 wire \soc/cpu/_04643_ ;
 wire \soc/cpu/_04644_ ;
 wire \soc/cpu/_04645_ ;
 wire \soc/cpu/_04646_ ;
 wire \soc/cpu/_04647_ ;
 wire \soc/cpu/_04648_ ;
 wire \soc/cpu/_04649_ ;
 wire \soc/cpu/_04650_ ;
 wire \soc/cpu/_04651_ ;
 wire \soc/cpu/_04652_ ;
 wire \soc/cpu/_04653_ ;
 wire \soc/cpu/_04654_ ;
 wire \soc/cpu/_04655_ ;
 wire \soc/cpu/_04656_ ;
 wire \soc/cpu/_04657_ ;
 wire \soc/cpu/_04658_ ;
 wire \soc/cpu/_04659_ ;
 wire \soc/cpu/_04660_ ;
 wire \soc/cpu/_04661_ ;
 wire \soc/cpu/_04662_ ;
 wire \soc/cpu/_04663_ ;
 wire \soc/cpu/_04664_ ;
 wire \soc/cpu/_04665_ ;
 wire \soc/cpu/_04666_ ;
 wire \soc/cpu/_04667_ ;
 wire \soc/cpu/_04668_ ;
 wire \soc/cpu/_04669_ ;
 wire net732;
 wire \soc/cpu/_04671_ ;
 wire \soc/cpu/_04672_ ;
 wire \soc/cpu/_04673_ ;
 wire \soc/cpu/_04674_ ;
 wire \soc/cpu/_04675_ ;
 wire \soc/cpu/_04676_ ;
 wire \soc/cpu/_04677_ ;
 wire \soc/cpu/_04678_ ;
 wire \soc/cpu/_04679_ ;
 wire \soc/cpu/_04680_ ;
 wire \soc/cpu/_04681_ ;
 wire \soc/cpu/_04682_ ;
 wire \soc/cpu/_04683_ ;
 wire \soc/cpu/_04684_ ;
 wire \soc/cpu/_04685_ ;
 wire \soc/cpu/_04686_ ;
 wire \soc/cpu/_04687_ ;
 wire \soc/cpu/_04688_ ;
 wire \soc/cpu/_04689_ ;
 wire \soc/cpu/_04690_ ;
 wire \soc/cpu/_04691_ ;
 wire \soc/cpu/_04692_ ;
 wire \soc/cpu/_04693_ ;
 wire \soc/cpu/_04694_ ;
 wire \soc/cpu/_04695_ ;
 wire \soc/cpu/_04696_ ;
 wire \soc/cpu/_04697_ ;
 wire \soc/cpu/_04698_ ;
 wire \soc/cpu/_04699_ ;
 wire \soc/cpu/_04700_ ;
 wire \soc/cpu/_04701_ ;
 wire \soc/cpu/_04702_ ;
 wire \soc/cpu/_04703_ ;
 wire \soc/cpu/_04704_ ;
 wire \soc/cpu/_04705_ ;
 wire \soc/cpu/_04706_ ;
 wire \soc/cpu/_04707_ ;
 wire \soc/cpu/_04708_ ;
 wire \soc/cpu/_04709_ ;
 wire \soc/cpu/_04710_ ;
 wire \soc/cpu/_04711_ ;
 wire \soc/cpu/_04712_ ;
 wire \soc/cpu/_04713_ ;
 wire \soc/cpu/_04714_ ;
 wire \soc/cpu/_04715_ ;
 wire \soc/cpu/_04716_ ;
 wire \soc/cpu/_04717_ ;
 wire \soc/cpu/_04718_ ;
 wire \soc/cpu/_04719_ ;
 wire \soc/cpu/_04720_ ;
 wire \soc/cpu/_04721_ ;
 wire \soc/cpu/_04722_ ;
 wire \soc/cpu/_04723_ ;
 wire \soc/cpu/_04724_ ;
 wire \soc/cpu/_04725_ ;
 wire \soc/cpu/_04726_ ;
 wire \soc/cpu/_04727_ ;
 wire \soc/cpu/_04728_ ;
 wire \soc/cpu/_04729_ ;
 wire \soc/cpu/_04730_ ;
 wire \soc/cpu/_04731_ ;
 wire \soc/cpu/_04732_ ;
 wire \soc/cpu/_04733_ ;
 wire \soc/cpu/_04734_ ;
 wire \soc/cpu/_04735_ ;
 wire \soc/cpu/_04736_ ;
 wire \soc/cpu/_04737_ ;
 wire \soc/cpu/_04738_ ;
 wire \soc/cpu/_04739_ ;
 wire \soc/cpu/_04740_ ;
 wire \soc/cpu/_04741_ ;
 wire \soc/cpu/_04742_ ;
 wire \soc/cpu/_04743_ ;
 wire \soc/cpu/_04744_ ;
 wire net731;
 wire net730;
 wire \soc/cpu/_04747_ ;
 wire net729;
 wire \soc/cpu/_04749_ ;
 wire net728;
 wire \soc/cpu/_04751_ ;
 wire \soc/cpu/_04752_ ;
 wire \soc/cpu/_04753_ ;
 wire \soc/cpu/_04754_ ;
 wire \soc/cpu/_04755_ ;
 wire \soc/cpu/_04756_ ;
 wire \soc/cpu/_04757_ ;
 wire \soc/cpu/_04758_ ;
 wire \soc/cpu/_04759_ ;
 wire net727;
 wire net726;
 wire \soc/cpu/_04762_ ;
 wire net725;
 wire \soc/cpu/_04764_ ;
 wire \soc/cpu/_04765_ ;
 wire \soc/cpu/_04766_ ;
 wire \soc/cpu/_04767_ ;
 wire \soc/cpu/_04768_ ;
 wire \soc/cpu/_04769_ ;
 wire \soc/cpu/_04770_ ;
 wire \soc/cpu/_04771_ ;
 wire \soc/cpu/_04772_ ;
 wire net724;
 wire net723;
 wire \soc/cpu/_04775_ ;
 wire net722;
 wire \soc/cpu/_04777_ ;
 wire \soc/cpu/_04778_ ;
 wire \soc/cpu/_04779_ ;
 wire \soc/cpu/_04780_ ;
 wire \soc/cpu/_04781_ ;
 wire \soc/cpu/_04782_ ;
 wire \soc/cpu/_04783_ ;
 wire \soc/cpu/_04784_ ;
 wire \soc/cpu/_04785_ ;
 wire \soc/cpu/_04786_ ;
 wire net721;
 wire \soc/cpu/_04788_ ;
 wire \soc/cpu/_04789_ ;
 wire \soc/cpu/_04790_ ;
 wire net720;
 wire \soc/cpu/_04792_ ;
 wire \soc/cpu/_04793_ ;
 wire net719;
 wire \soc/cpu/_04795_ ;
 wire \soc/cpu/_04796_ ;
 wire \soc/cpu/_04797_ ;
 wire \soc/cpu/_04798_ ;
 wire \soc/cpu/_04799_ ;
 wire \soc/cpu/_04800_ ;
 wire \soc/cpu/_04801_ ;
 wire \soc/cpu/_04802_ ;
 wire \soc/cpu/_04803_ ;
 wire \soc/cpu/_04804_ ;
 wire \soc/cpu/_04805_ ;
 wire \soc/cpu/_04806_ ;
 wire \soc/cpu/_04807_ ;
 wire \soc/cpu/_04808_ ;
 wire \soc/cpu/_04809_ ;
 wire net718;
 wire \soc/cpu/_04811_ ;
 wire \soc/cpu/_04812_ ;
 wire net717;
 wire net716;
 wire \soc/cpu/_04815_ ;
 wire \soc/cpu/_04816_ ;
 wire \soc/cpu/_04817_ ;
 wire \soc/cpu/_04818_ ;
 wire \soc/cpu/_04819_ ;
 wire \soc/cpu/_04820_ ;
 wire \soc/cpu/_04821_ ;
 wire \soc/cpu/_04822_ ;
 wire \soc/cpu/_04823_ ;
 wire \soc/cpu/_04824_ ;
 wire \soc/cpu/_04825_ ;
 wire \soc/cpu/_04826_ ;
 wire \soc/cpu/_04827_ ;
 wire \soc/cpu/_04828_ ;
 wire \soc/cpu/_04829_ ;
 wire \soc/cpu/_04830_ ;
 wire net715;
 wire \soc/cpu/_04832_ ;
 wire \soc/cpu/_04833_ ;
 wire \soc/cpu/_04834_ ;
 wire \soc/cpu/_04835_ ;
 wire net714;
 wire net713;
 wire \soc/cpu/_04838_ ;
 wire \soc/cpu/_04839_ ;
 wire \soc/cpu/_04840_ ;
 wire \soc/cpu/_04841_ ;
 wire \soc/cpu/_04842_ ;
 wire \soc/cpu/_04843_ ;
 wire \soc/cpu/_04844_ ;
 wire \soc/cpu/_04845_ ;
 wire \soc/cpu/_04846_ ;
 wire \soc/cpu/_04847_ ;
 wire \soc/cpu/_04848_ ;
 wire \soc/cpu/_04849_ ;
 wire \soc/cpu/_04850_ ;
 wire \soc/cpu/_04851_ ;
 wire \soc/cpu/_04852_ ;
 wire \soc/cpu/_04853_ ;
 wire \soc/cpu/_04854_ ;
 wire \soc/cpu/_04855_ ;
 wire \soc/cpu/_04856_ ;
 wire \soc/cpu/_04857_ ;
 wire \soc/cpu/_04858_ ;
 wire \soc/cpu/_04859_ ;
 wire \soc/cpu/_04860_ ;
 wire \soc/cpu/_04861_ ;
 wire \soc/cpu/_04862_ ;
 wire \soc/cpu/_04863_ ;
 wire \soc/cpu/_04864_ ;
 wire \soc/cpu/_04865_ ;
 wire \soc/cpu/_04866_ ;
 wire \soc/cpu/_04867_ ;
 wire \soc/cpu/_04868_ ;
 wire net458;
 wire \soc/cpu/alu_out[0] ;
 wire \soc/cpu/alu_out[10] ;
 wire \soc/cpu/alu_out[11] ;
 wire \soc/cpu/alu_out[12] ;
 wire \soc/cpu/alu_out[13] ;
 wire \soc/cpu/alu_out[14] ;
 wire \soc/cpu/alu_out[15] ;
 wire \soc/cpu/alu_out[16] ;
 wire \soc/cpu/alu_out[17] ;
 wire \soc/cpu/alu_out[18] ;
 wire \soc/cpu/alu_out[19] ;
 wire \soc/cpu/alu_out[1] ;
 wire \soc/cpu/alu_out[20] ;
 wire \soc/cpu/alu_out[21] ;
 wire \soc/cpu/alu_out[22] ;
 wire \soc/cpu/alu_out[23] ;
 wire \soc/cpu/alu_out[24] ;
 wire \soc/cpu/alu_out[25] ;
 wire \soc/cpu/alu_out[26] ;
 wire \soc/cpu/alu_out[27] ;
 wire \soc/cpu/alu_out[28] ;
 wire \soc/cpu/alu_out[29] ;
 wire \soc/cpu/alu_out[2] ;
 wire \soc/cpu/alu_out[30] ;
 wire \soc/cpu/alu_out[31] ;
 wire \soc/cpu/alu_out[3] ;
 wire \soc/cpu/alu_out[4] ;
 wire \soc/cpu/alu_out[5] ;
 wire \soc/cpu/alu_out[6] ;
 wire \soc/cpu/alu_out[7] ;
 wire \soc/cpu/alu_out[8] ;
 wire \soc/cpu/alu_out[9] ;
 wire \soc/cpu/alu_out_q[0] ;
 wire \soc/cpu/alu_out_q[10] ;
 wire \soc/cpu/alu_out_q[11] ;
 wire \soc/cpu/alu_out_q[12] ;
 wire \soc/cpu/alu_out_q[13] ;
 wire \soc/cpu/alu_out_q[14] ;
 wire \soc/cpu/alu_out_q[15] ;
 wire \soc/cpu/alu_out_q[16] ;
 wire \soc/cpu/alu_out_q[17] ;
 wire \soc/cpu/alu_out_q[18] ;
 wire \soc/cpu/alu_out_q[19] ;
 wire \soc/cpu/alu_out_q[1] ;
 wire \soc/cpu/alu_out_q[20] ;
 wire \soc/cpu/alu_out_q[21] ;
 wire \soc/cpu/alu_out_q[22] ;
 wire \soc/cpu/alu_out_q[23] ;
 wire \soc/cpu/alu_out_q[24] ;
 wire \soc/cpu/alu_out_q[25] ;
 wire \soc/cpu/alu_out_q[26] ;
 wire \soc/cpu/alu_out_q[27] ;
 wire \soc/cpu/alu_out_q[28] ;
 wire \soc/cpu/alu_out_q[29] ;
 wire \soc/cpu/alu_out_q[2] ;
 wire \soc/cpu/alu_out_q[30] ;
 wire \soc/cpu/alu_out_q[31] ;
 wire \soc/cpu/alu_out_q[3] ;
 wire \soc/cpu/alu_out_q[4] ;
 wire \soc/cpu/alu_out_q[5] ;
 wire \soc/cpu/alu_out_q[6] ;
 wire \soc/cpu/alu_out_q[7] ;
 wire \soc/cpu/alu_out_q[8] ;
 wire \soc/cpu/alu_out_q[9] ;
 wire \soc/cpu/clear_prefetched_high_word ;
 wire \soc/cpu/clear_prefetched_high_word_q ;
 wire \soc/cpu/compressed_instr ;
 wire \soc/cpu/count_cycle[0] ;
 wire \soc/cpu/count_cycle[10] ;
 wire \soc/cpu/count_cycle[11] ;
 wire \soc/cpu/count_cycle[12] ;
 wire \soc/cpu/count_cycle[13] ;
 wire \soc/cpu/count_cycle[14] ;
 wire \soc/cpu/count_cycle[15] ;
 wire \soc/cpu/count_cycle[16] ;
 wire \soc/cpu/count_cycle[17] ;
 wire \soc/cpu/count_cycle[18] ;
 wire \soc/cpu/count_cycle[19] ;
 wire \soc/cpu/count_cycle[1] ;
 wire \soc/cpu/count_cycle[20] ;
 wire \soc/cpu/count_cycle[21] ;
 wire \soc/cpu/count_cycle[22] ;
 wire \soc/cpu/count_cycle[23] ;
 wire \soc/cpu/count_cycle[24] ;
 wire \soc/cpu/count_cycle[25] ;
 wire \soc/cpu/count_cycle[26] ;
 wire \soc/cpu/count_cycle[27] ;
 wire \soc/cpu/count_cycle[28] ;
 wire \soc/cpu/count_cycle[29] ;
 wire \soc/cpu/count_cycle[2] ;
 wire \soc/cpu/count_cycle[30] ;
 wire \soc/cpu/count_cycle[31] ;
 wire \soc/cpu/count_cycle[32] ;
 wire \soc/cpu/count_cycle[33] ;
 wire \soc/cpu/count_cycle[34] ;
 wire \soc/cpu/count_cycle[35] ;
 wire \soc/cpu/count_cycle[36] ;
 wire \soc/cpu/count_cycle[37] ;
 wire \soc/cpu/count_cycle[38] ;
 wire \soc/cpu/count_cycle[39] ;
 wire \soc/cpu/count_cycle[3] ;
 wire \soc/cpu/count_cycle[40] ;
 wire \soc/cpu/count_cycle[41] ;
 wire \soc/cpu/count_cycle[42] ;
 wire \soc/cpu/count_cycle[43] ;
 wire \soc/cpu/count_cycle[44] ;
 wire \soc/cpu/count_cycle[45] ;
 wire \soc/cpu/count_cycle[46] ;
 wire \soc/cpu/count_cycle[47] ;
 wire \soc/cpu/count_cycle[48] ;
 wire \soc/cpu/count_cycle[49] ;
 wire \soc/cpu/count_cycle[4] ;
 wire \soc/cpu/count_cycle[50] ;
 wire \soc/cpu/count_cycle[51] ;
 wire \soc/cpu/count_cycle[52] ;
 wire \soc/cpu/count_cycle[53] ;
 wire \soc/cpu/count_cycle[54] ;
 wire \soc/cpu/count_cycle[55] ;
 wire \soc/cpu/count_cycle[56] ;
 wire \soc/cpu/count_cycle[57] ;
 wire \soc/cpu/count_cycle[58] ;
 wire \soc/cpu/count_cycle[59] ;
 wire \soc/cpu/count_cycle[5] ;
 wire \soc/cpu/count_cycle[60] ;
 wire \soc/cpu/count_cycle[61] ;
 wire \soc/cpu/count_cycle[62] ;
 wire \soc/cpu/count_cycle[63] ;
 wire \soc/cpu/count_cycle[6] ;
 wire \soc/cpu/count_cycle[7] ;
 wire \soc/cpu/count_cycle[8] ;
 wire \soc/cpu/count_cycle[9] ;
 wire \soc/cpu/count_instr[0] ;
 wire \soc/cpu/count_instr[10] ;
 wire \soc/cpu/count_instr[11] ;
 wire \soc/cpu/count_instr[12] ;
 wire \soc/cpu/count_instr[13] ;
 wire \soc/cpu/count_instr[14] ;
 wire \soc/cpu/count_instr[15] ;
 wire \soc/cpu/count_instr[16] ;
 wire \soc/cpu/count_instr[17] ;
 wire \soc/cpu/count_instr[18] ;
 wire \soc/cpu/count_instr[19] ;
 wire \soc/cpu/count_instr[1] ;
 wire \soc/cpu/count_instr[20] ;
 wire \soc/cpu/count_instr[21] ;
 wire \soc/cpu/count_instr[22] ;
 wire \soc/cpu/count_instr[23] ;
 wire \soc/cpu/count_instr[24] ;
 wire \soc/cpu/count_instr[25] ;
 wire \soc/cpu/count_instr[26] ;
 wire \soc/cpu/count_instr[27] ;
 wire \soc/cpu/count_instr[28] ;
 wire \soc/cpu/count_instr[29] ;
 wire \soc/cpu/count_instr[2] ;
 wire \soc/cpu/count_instr[30] ;
 wire \soc/cpu/count_instr[31] ;
 wire \soc/cpu/count_instr[32] ;
 wire \soc/cpu/count_instr[33] ;
 wire \soc/cpu/count_instr[34] ;
 wire \soc/cpu/count_instr[35] ;
 wire \soc/cpu/count_instr[36] ;
 wire \soc/cpu/count_instr[37] ;
 wire \soc/cpu/count_instr[38] ;
 wire \soc/cpu/count_instr[39] ;
 wire \soc/cpu/count_instr[3] ;
 wire \soc/cpu/count_instr[40] ;
 wire \soc/cpu/count_instr[41] ;
 wire \soc/cpu/count_instr[42] ;
 wire \soc/cpu/count_instr[43] ;
 wire \soc/cpu/count_instr[44] ;
 wire \soc/cpu/count_instr[45] ;
 wire \soc/cpu/count_instr[46] ;
 wire \soc/cpu/count_instr[47] ;
 wire \soc/cpu/count_instr[48] ;
 wire \soc/cpu/count_instr[49] ;
 wire \soc/cpu/count_instr[4] ;
 wire \soc/cpu/count_instr[50] ;
 wire \soc/cpu/count_instr[51] ;
 wire \soc/cpu/count_instr[52] ;
 wire \soc/cpu/count_instr[53] ;
 wire \soc/cpu/count_instr[54] ;
 wire \soc/cpu/count_instr[55] ;
 wire \soc/cpu/count_instr[56] ;
 wire \soc/cpu/count_instr[57] ;
 wire \soc/cpu/count_instr[58] ;
 wire \soc/cpu/count_instr[59] ;
 wire \soc/cpu/count_instr[5] ;
 wire \soc/cpu/count_instr[60] ;
 wire \soc/cpu/count_instr[61] ;
 wire \soc/cpu/count_instr[62] ;
 wire \soc/cpu/count_instr[63] ;
 wire \soc/cpu/count_instr[6] ;
 wire \soc/cpu/count_instr[7] ;
 wire \soc/cpu/count_instr[8] ;
 wire \soc/cpu/count_instr[9] ;
 wire \soc/cpu/cpu_state[0] ;
 wire \soc/cpu/cpu_state[1] ;
 wire \soc/cpu/cpu_state[2] ;
 wire \soc/cpu/cpu_state[3] ;
 wire \soc/cpu/cpu_state[4] ;
 wire \soc/cpu/cpu_state[5] ;
 wire \soc/cpu/cpu_state[6] ;
 wire \soc/cpu/cpuregs_raddr1[0] ;
 wire \soc/cpu/cpuregs_raddr1[1] ;
 wire \soc/cpu/cpuregs_raddr1[2] ;
 wire \soc/cpu/cpuregs_raddr1[3] ;
 wire \soc/cpu/cpuregs_raddr1[4] ;
 wire \soc/cpu/cpuregs_raddr2[0] ;
 wire \soc/cpu/cpuregs_raddr2[1] ;
 wire \soc/cpu/cpuregs_raddr2[2] ;
 wire \soc/cpu/cpuregs_raddr2[3] ;
 wire \soc/cpu/cpuregs_raddr2[4] ;
 wire \soc/cpu/cpuregs_rdata1[0] ;
 wire \soc/cpu/cpuregs_rdata1[10] ;
 wire \soc/cpu/cpuregs_rdata1[11] ;
 wire \soc/cpu/cpuregs_rdata1[12] ;
 wire \soc/cpu/cpuregs_rdata1[13] ;
 wire \soc/cpu/cpuregs_rdata1[14] ;
 wire \soc/cpu/cpuregs_rdata1[15] ;
 wire \soc/cpu/cpuregs_rdata1[16] ;
 wire \soc/cpu/cpuregs_rdata1[17] ;
 wire \soc/cpu/cpuregs_rdata1[18] ;
 wire \soc/cpu/cpuregs_rdata1[19] ;
 wire \soc/cpu/cpuregs_rdata1[1] ;
 wire \soc/cpu/cpuregs_rdata1[20] ;
 wire \soc/cpu/cpuregs_rdata1[21] ;
 wire \soc/cpu/cpuregs_rdata1[22] ;
 wire \soc/cpu/cpuregs_rdata1[23] ;
 wire \soc/cpu/cpuregs_rdata1[24] ;
 wire \soc/cpu/cpuregs_rdata1[25] ;
 wire \soc/cpu/cpuregs_rdata1[26] ;
 wire \soc/cpu/cpuregs_rdata1[27] ;
 wire \soc/cpu/cpuregs_rdata1[28] ;
 wire \soc/cpu/cpuregs_rdata1[29] ;
 wire \soc/cpu/cpuregs_rdata1[2] ;
 wire \soc/cpu/cpuregs_rdata1[30] ;
 wire \soc/cpu/cpuregs_rdata1[31] ;
 wire \soc/cpu/cpuregs_rdata1[3] ;
 wire \soc/cpu/cpuregs_rdata1[4] ;
 wire \soc/cpu/cpuregs_rdata1[5] ;
 wire \soc/cpu/cpuregs_rdata1[6] ;
 wire \soc/cpu/cpuregs_rdata1[7] ;
 wire \soc/cpu/cpuregs_rdata1[8] ;
 wire \soc/cpu/cpuregs_rdata1[9] ;
 wire \soc/cpu/cpuregs_rdata2[0] ;
 wire \soc/cpu/cpuregs_rdata2[10] ;
 wire \soc/cpu/cpuregs_rdata2[11] ;
 wire \soc/cpu/cpuregs_rdata2[12] ;
 wire \soc/cpu/cpuregs_rdata2[13] ;
 wire \soc/cpu/cpuregs_rdata2[14] ;
 wire \soc/cpu/cpuregs_rdata2[15] ;
 wire \soc/cpu/cpuregs_rdata2[16] ;
 wire \soc/cpu/cpuregs_rdata2[17] ;
 wire \soc/cpu/cpuregs_rdata2[18] ;
 wire \soc/cpu/cpuregs_rdata2[19] ;
 wire \soc/cpu/cpuregs_rdata2[1] ;
 wire \soc/cpu/cpuregs_rdata2[20] ;
 wire \soc/cpu/cpuregs_rdata2[21] ;
 wire \soc/cpu/cpuregs_rdata2[22] ;
 wire \soc/cpu/cpuregs_rdata2[23] ;
 wire \soc/cpu/cpuregs_rdata2[24] ;
 wire \soc/cpu/cpuregs_rdata2[25] ;
 wire \soc/cpu/cpuregs_rdata2[26] ;
 wire \soc/cpu/cpuregs_rdata2[27] ;
 wire \soc/cpu/cpuregs_rdata2[28] ;
 wire \soc/cpu/cpuregs_rdata2[29] ;
 wire \soc/cpu/cpuregs_rdata2[2] ;
 wire \soc/cpu/cpuregs_rdata2[30] ;
 wire \soc/cpu/cpuregs_rdata2[31] ;
 wire \soc/cpu/cpuregs_rdata2[3] ;
 wire \soc/cpu/cpuregs_rdata2[4] ;
 wire \soc/cpu/cpuregs_rdata2[5] ;
 wire \soc/cpu/cpuregs_rdata2[6] ;
 wire \soc/cpu/cpuregs_rdata2[7] ;
 wire \soc/cpu/cpuregs_rdata2[8] ;
 wire \soc/cpu/cpuregs_rdata2[9] ;
 wire \soc/cpu/cpuregs_waddr[0] ;
 wire \soc/cpu/cpuregs_waddr[1] ;
 wire \soc/cpu/cpuregs_waddr[2] ;
 wire \soc/cpu/cpuregs_waddr[3] ;
 wire \soc/cpu/cpuregs_waddr[4] ;
 wire \soc/cpu/cpuregs_wrdata[0] ;
 wire \soc/cpu/cpuregs_wrdata[10] ;
 wire \soc/cpu/cpuregs_wrdata[11] ;
 wire \soc/cpu/cpuregs_wrdata[12] ;
 wire \soc/cpu/cpuregs_wrdata[13] ;
 wire \soc/cpu/cpuregs_wrdata[14] ;
 wire \soc/cpu/cpuregs_wrdata[15] ;
 wire \soc/cpu/cpuregs_wrdata[16] ;
 wire \soc/cpu/cpuregs_wrdata[17] ;
 wire \soc/cpu/cpuregs_wrdata[18] ;
 wire \soc/cpu/cpuregs_wrdata[19] ;
 wire \soc/cpu/cpuregs_wrdata[1] ;
 wire \soc/cpu/cpuregs_wrdata[20] ;
 wire \soc/cpu/cpuregs_wrdata[21] ;
 wire \soc/cpu/cpuregs_wrdata[22] ;
 wire \soc/cpu/cpuregs_wrdata[23] ;
 wire \soc/cpu/cpuregs_wrdata[24] ;
 wire \soc/cpu/cpuregs_wrdata[25] ;
 wire \soc/cpu/cpuregs_wrdata[26] ;
 wire \soc/cpu/cpuregs_wrdata[27] ;
 wire \soc/cpu/cpuregs_wrdata[28] ;
 wire \soc/cpu/cpuregs_wrdata[29] ;
 wire \soc/cpu/cpuregs_wrdata[2] ;
 wire \soc/cpu/cpuregs_wrdata[30] ;
 wire \soc/cpu/cpuregs_wrdata[31] ;
 wire \soc/cpu/cpuregs_wrdata[3] ;
 wire \soc/cpu/cpuregs_wrdata[4] ;
 wire \soc/cpu/cpuregs_wrdata[5] ;
 wire \soc/cpu/cpuregs_wrdata[6] ;
 wire \soc/cpu/cpuregs_wrdata[7] ;
 wire \soc/cpu/cpuregs_wrdata[8] ;
 wire \soc/cpu/cpuregs_wrdata[9] ;
 wire \soc/cpu/decoded_imm[0] ;
 wire \soc/cpu/decoded_imm[10] ;
 wire \soc/cpu/decoded_imm[11] ;
 wire \soc/cpu/decoded_imm[12] ;
 wire \soc/cpu/decoded_imm[13] ;
 wire \soc/cpu/decoded_imm[14] ;
 wire \soc/cpu/decoded_imm[15] ;
 wire \soc/cpu/decoded_imm[16] ;
 wire \soc/cpu/decoded_imm[17] ;
 wire \soc/cpu/decoded_imm[18] ;
 wire \soc/cpu/decoded_imm[19] ;
 wire \soc/cpu/decoded_imm[1] ;
 wire \soc/cpu/decoded_imm[20] ;
 wire \soc/cpu/decoded_imm[21] ;
 wire \soc/cpu/decoded_imm[22] ;
 wire \soc/cpu/decoded_imm[23] ;
 wire \soc/cpu/decoded_imm[24] ;
 wire \soc/cpu/decoded_imm[25] ;
 wire \soc/cpu/decoded_imm[26] ;
 wire \soc/cpu/decoded_imm[27] ;
 wire \soc/cpu/decoded_imm[28] ;
 wire \soc/cpu/decoded_imm[29] ;
 wire \soc/cpu/decoded_imm[2] ;
 wire \soc/cpu/decoded_imm[30] ;
 wire \soc/cpu/decoded_imm[31] ;
 wire \soc/cpu/decoded_imm[3] ;
 wire \soc/cpu/decoded_imm[4] ;
 wire \soc/cpu/decoded_imm[5] ;
 wire \soc/cpu/decoded_imm[6] ;
 wire \soc/cpu/decoded_imm[7] ;
 wire \soc/cpu/decoded_imm[8] ;
 wire \soc/cpu/decoded_imm[9] ;
 wire \soc/cpu/decoded_imm_j[10] ;
 wire \soc/cpu/decoded_imm_j[11] ;
 wire \soc/cpu/decoded_imm_j[12] ;
 wire \soc/cpu/decoded_imm_j[13] ;
 wire \soc/cpu/decoded_imm_j[14] ;
 wire \soc/cpu/decoded_imm_j[15] ;
 wire \soc/cpu/decoded_imm_j[16] ;
 wire \soc/cpu/decoded_imm_j[17] ;
 wire \soc/cpu/decoded_imm_j[18] ;
 wire \soc/cpu/decoded_imm_j[19] ;
 wire \soc/cpu/decoded_imm_j[1] ;
 wire \soc/cpu/decoded_imm_j[20] ;
 wire \soc/cpu/decoded_imm_j[2] ;
 wire \soc/cpu/decoded_imm_j[3] ;
 wire \soc/cpu/decoded_imm_j[4] ;
 wire \soc/cpu/decoded_imm_j[5] ;
 wire \soc/cpu/decoded_imm_j[6] ;
 wire \soc/cpu/decoded_imm_j[7] ;
 wire \soc/cpu/decoded_imm_j[8] ;
 wire \soc/cpu/decoded_imm_j[9] ;
 wire \soc/cpu/decoded_rd[0] ;
 wire \soc/cpu/decoded_rd[1] ;
 wire \soc/cpu/decoded_rd[2] ;
 wire \soc/cpu/decoded_rd[3] ;
 wire \soc/cpu/decoded_rd[4] ;
 wire \soc/cpu/decoder_pseudo_trigger ;
 wire \soc/cpu/decoder_trigger ;
 wire \soc/cpu/do_waitirq ;
 wire \soc/cpu/instr_add ;
 wire \soc/cpu/instr_addi ;
 wire \soc/cpu/instr_and ;
 wire \soc/cpu/instr_andi ;
 wire \soc/cpu/instr_auipc ;
 wire \soc/cpu/instr_beq ;
 wire \soc/cpu/instr_bge ;
 wire \soc/cpu/instr_bgeu ;
 wire \soc/cpu/instr_blt ;
 wire \soc/cpu/instr_bltu ;
 wire \soc/cpu/instr_bne ;
 wire \soc/cpu/instr_fence ;
 wire \soc/cpu/instr_jal ;
 wire \soc/cpu/instr_jalr ;
 wire \soc/cpu/instr_lb ;
 wire \soc/cpu/instr_lbu ;
 wire \soc/cpu/instr_lh ;
 wire \soc/cpu/instr_lhu ;
 wire \soc/cpu/instr_lui ;
 wire \soc/cpu/instr_lw ;
 wire \soc/cpu/instr_maskirq ;
 wire \soc/cpu/instr_or ;
 wire \soc/cpu/instr_ori ;
 wire \soc/cpu/instr_rdcycle ;
 wire \soc/cpu/instr_rdcycleh ;
 wire \soc/cpu/instr_rdinstr ;
 wire \soc/cpu/instr_rdinstrh ;
 wire \soc/cpu/instr_retirq ;
 wire \soc/cpu/instr_sb ;
 wire \soc/cpu/instr_sh ;
 wire \soc/cpu/instr_sll ;
 wire \soc/cpu/instr_slli ;
 wire \soc/cpu/instr_slt ;
 wire \soc/cpu/instr_slti ;
 wire \soc/cpu/instr_sltiu ;
 wire \soc/cpu/instr_sltu ;
 wire \soc/cpu/instr_sra ;
 wire \soc/cpu/instr_srai ;
 wire \soc/cpu/instr_srl ;
 wire \soc/cpu/instr_srli ;
 wire \soc/cpu/instr_sub ;
 wire \soc/cpu/instr_sw ;
 wire \soc/cpu/instr_timer ;
 wire \soc/cpu/instr_waitirq ;
 wire \soc/cpu/instr_xor ;
 wire \soc/cpu/instr_xori ;
 wire \soc/cpu/irq_active ;
 wire \soc/cpu/irq_delay ;
 wire \soc/cpu/irq_mask[0] ;
 wire \soc/cpu/irq_mask[10] ;
 wire \soc/cpu/irq_mask[11] ;
 wire \soc/cpu/irq_mask[12] ;
 wire \soc/cpu/irq_mask[13] ;
 wire \soc/cpu/irq_mask[14] ;
 wire \soc/cpu/irq_mask[15] ;
 wire \soc/cpu/irq_mask[16] ;
 wire \soc/cpu/irq_mask[17] ;
 wire \soc/cpu/irq_mask[18] ;
 wire \soc/cpu/irq_mask[19] ;
 wire \soc/cpu/irq_mask[1] ;
 wire \soc/cpu/irq_mask[20] ;
 wire \soc/cpu/irq_mask[21] ;
 wire \soc/cpu/irq_mask[22] ;
 wire \soc/cpu/irq_mask[23] ;
 wire \soc/cpu/irq_mask[24] ;
 wire \soc/cpu/irq_mask[25] ;
 wire \soc/cpu/irq_mask[26] ;
 wire \soc/cpu/irq_mask[27] ;
 wire \soc/cpu/irq_mask[28] ;
 wire \soc/cpu/irq_mask[29] ;
 wire \soc/cpu/irq_mask[2] ;
 wire \soc/cpu/irq_mask[30] ;
 wire \soc/cpu/irq_mask[31] ;
 wire \soc/cpu/irq_mask[3] ;
 wire \soc/cpu/irq_mask[4] ;
 wire \soc/cpu/irq_mask[5] ;
 wire \soc/cpu/irq_mask[6] ;
 wire \soc/cpu/irq_mask[7] ;
 wire \soc/cpu/irq_mask[8] ;
 wire \soc/cpu/irq_mask[9] ;
 wire \soc/cpu/irq_pending[0] ;
 wire \soc/cpu/irq_pending[10] ;
 wire \soc/cpu/irq_pending[11] ;
 wire \soc/cpu/irq_pending[12] ;
 wire \soc/cpu/irq_pending[13] ;
 wire \soc/cpu/irq_pending[14] ;
 wire \soc/cpu/irq_pending[15] ;
 wire \soc/cpu/irq_pending[16] ;
 wire \soc/cpu/irq_pending[17] ;
 wire \soc/cpu/irq_pending[18] ;
 wire \soc/cpu/irq_pending[19] ;
 wire \soc/cpu/irq_pending[1] ;
 wire \soc/cpu/irq_pending[20] ;
 wire \soc/cpu/irq_pending[21] ;
 wire \soc/cpu/irq_pending[22] ;
 wire \soc/cpu/irq_pending[23] ;
 wire \soc/cpu/irq_pending[24] ;
 wire \soc/cpu/irq_pending[25] ;
 wire \soc/cpu/irq_pending[26] ;
 wire \soc/cpu/irq_pending[27] ;
 wire \soc/cpu/irq_pending[28] ;
 wire \soc/cpu/irq_pending[29] ;
 wire \soc/cpu/irq_pending[2] ;
 wire \soc/cpu/irq_pending[30] ;
 wire \soc/cpu/irq_pending[31] ;
 wire \soc/cpu/irq_pending[3] ;
 wire \soc/cpu/irq_pending[4] ;
 wire \soc/cpu/irq_pending[5] ;
 wire \soc/cpu/irq_pending[6] ;
 wire \soc/cpu/irq_pending[7] ;
 wire \soc/cpu/irq_pending[8] ;
 wire \soc/cpu/irq_pending[9] ;
 wire \soc/cpu/irq_state[0] ;
 wire \soc/cpu/irq_state[1] ;
 wire \soc/cpu/is_alu_reg_imm ;
 wire \soc/cpu/is_alu_reg_reg ;
 wire \soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ;
 wire \soc/cpu/is_compare ;
 wire \soc/cpu/is_jalr_addi_slti_sltiu_xori_ori_andi ;
 wire \soc/cpu/is_lb_lh_lw_lbu_lhu ;
 wire \soc/cpu/is_lui_auipc_jal ;
 wire \soc/cpu/is_sb_sh_sw ;
 wire \soc/cpu/is_sll_srl_sra ;
 wire \soc/cpu/is_slli_srli_srai ;
 wire \soc/cpu/is_slti_blt_slt ;
 wire \soc/cpu/is_sltiu_bltu_sltu ;
 wire \soc/cpu/last_mem_valid ;
 wire \soc/cpu/latched_branch ;
 wire \soc/cpu/latched_compr ;
 wire \soc/cpu/latched_is_lb ;
 wire \soc/cpu/latched_is_lh ;
 wire \soc/cpu/latched_stalu ;
 wire \soc/cpu/latched_store ;
 wire \soc/cpu/mem_16bit_buffer[0] ;
 wire \soc/cpu/mem_16bit_buffer[10] ;
 wire \soc/cpu/mem_16bit_buffer[11] ;
 wire \soc/cpu/mem_16bit_buffer[12] ;
 wire \soc/cpu/mem_16bit_buffer[13] ;
 wire \soc/cpu/mem_16bit_buffer[14] ;
 wire \soc/cpu/mem_16bit_buffer[15] ;
 wire \soc/cpu/mem_16bit_buffer[1] ;
 wire \soc/cpu/mem_16bit_buffer[2] ;
 wire \soc/cpu/mem_16bit_buffer[3] ;
 wire \soc/cpu/mem_16bit_buffer[4] ;
 wire \soc/cpu/mem_16bit_buffer[5] ;
 wire \soc/cpu/mem_16bit_buffer[6] ;
 wire \soc/cpu/mem_16bit_buffer[7] ;
 wire \soc/cpu/mem_16bit_buffer[8] ;
 wire \soc/cpu/mem_16bit_buffer[9] ;
 wire \soc/cpu/mem_do_prefetch ;
 wire \soc/cpu/mem_do_rdata ;
 wire \soc/cpu/mem_do_rinst ;
 wire \soc/cpu/mem_do_wdata ;
 wire net710;
 wire net709;
 wire \soc/cpu/mem_la_firstword_reg ;
 wire \soc/cpu/mem_la_read ;
 wire \soc/cpu/mem_la_secondword ;
 wire \soc/cpu/mem_rdata_q[0] ;
 wire \soc/cpu/mem_rdata_q[10] ;
 wire \soc/cpu/mem_rdata_q[11] ;
 wire \soc/cpu/mem_rdata_q[12] ;
 wire \soc/cpu/mem_rdata_q[13] ;
 wire \soc/cpu/mem_rdata_q[14] ;
 wire \soc/cpu/mem_rdata_q[15] ;
 wire \soc/cpu/mem_rdata_q[16] ;
 wire \soc/cpu/mem_rdata_q[17] ;
 wire \soc/cpu/mem_rdata_q[18] ;
 wire \soc/cpu/mem_rdata_q[19] ;
 wire \soc/cpu/mem_rdata_q[1] ;
 wire \soc/cpu/mem_rdata_q[20] ;
 wire \soc/cpu/mem_rdata_q[21] ;
 wire \soc/cpu/mem_rdata_q[22] ;
 wire \soc/cpu/mem_rdata_q[23] ;
 wire \soc/cpu/mem_rdata_q[24] ;
 wire \soc/cpu/mem_rdata_q[25] ;
 wire \soc/cpu/mem_rdata_q[26] ;
 wire \soc/cpu/mem_rdata_q[27] ;
 wire \soc/cpu/mem_rdata_q[28] ;
 wire \soc/cpu/mem_rdata_q[29] ;
 wire \soc/cpu/mem_rdata_q[2] ;
 wire \soc/cpu/mem_rdata_q[30] ;
 wire \soc/cpu/mem_rdata_q[31] ;
 wire \soc/cpu/mem_rdata_q[3] ;
 wire \soc/cpu/mem_rdata_q[4] ;
 wire \soc/cpu/mem_rdata_q[5] ;
 wire \soc/cpu/mem_rdata_q[6] ;
 wire \soc/cpu/mem_rdata_q[7] ;
 wire \soc/cpu/mem_rdata_q[8] ;
 wire \soc/cpu/mem_rdata_q[9] ;
 wire \soc/cpu/mem_state[0] ;
 wire \soc/cpu/mem_state[1] ;
 wire \soc/cpu/mem_wordsize[0] ;
 wire \soc/cpu/mem_wordsize[1] ;
 wire \soc/cpu/mem_wordsize[2] ;
 wire net708;
 wire net698;
 wire net697;
 wire net696;
 wire net695;
 wire net694;
 wire net693;
 wire net692;
 wire net691;
 wire net690;
 wire net689;
 wire net707;
 wire net688;
 wire net687;
 wire net686;
 wire net685;
 wire net684;
 wire net683;
 wire net682;
 wire net681;
 wire net680;
 wire net679;
 wire net706;
 wire net678;
 wire net677;
 wire net705;
 wire net704;
 wire net703;
 wire net702;
 wire net701;
 wire net700;
 wire net699;
 wire net676;
 wire net675;
 wire net674;
 wire net673;
 wire net672;
 wire net671;
 wire net670;
 wire net669;
 wire net668;
 wire \soc/cpu/prefetched_high_word ;
 wire \soc/cpu/reg_next_pc[0] ;
 wire \soc/cpu/reg_next_pc[10] ;
 wire \soc/cpu/reg_next_pc[11] ;
 wire \soc/cpu/reg_next_pc[12] ;
 wire \soc/cpu/reg_next_pc[13] ;
 wire \soc/cpu/reg_next_pc[14] ;
 wire \soc/cpu/reg_next_pc[15] ;
 wire \soc/cpu/reg_next_pc[16] ;
 wire \soc/cpu/reg_next_pc[17] ;
 wire \soc/cpu/reg_next_pc[18] ;
 wire \soc/cpu/reg_next_pc[19] ;
 wire \soc/cpu/reg_next_pc[1] ;
 wire \soc/cpu/reg_next_pc[20] ;
 wire \soc/cpu/reg_next_pc[21] ;
 wire \soc/cpu/reg_next_pc[22] ;
 wire \soc/cpu/reg_next_pc[23] ;
 wire \soc/cpu/reg_next_pc[24] ;
 wire \soc/cpu/reg_next_pc[25] ;
 wire \soc/cpu/reg_next_pc[26] ;
 wire \soc/cpu/reg_next_pc[27] ;
 wire \soc/cpu/reg_next_pc[28] ;
 wire \soc/cpu/reg_next_pc[29] ;
 wire \soc/cpu/reg_next_pc[2] ;
 wire \soc/cpu/reg_next_pc[30] ;
 wire \soc/cpu/reg_next_pc[31] ;
 wire \soc/cpu/reg_next_pc[3] ;
 wire \soc/cpu/reg_next_pc[4] ;
 wire \soc/cpu/reg_next_pc[5] ;
 wire \soc/cpu/reg_next_pc[6] ;
 wire \soc/cpu/reg_next_pc[7] ;
 wire \soc/cpu/reg_next_pc[8] ;
 wire \soc/cpu/reg_next_pc[9] ;
 wire \soc/cpu/reg_out[0] ;
 wire \soc/cpu/reg_out[10] ;
 wire \soc/cpu/reg_out[11] ;
 wire \soc/cpu/reg_out[12] ;
 wire \soc/cpu/reg_out[13] ;
 wire \soc/cpu/reg_out[14] ;
 wire \soc/cpu/reg_out[15] ;
 wire \soc/cpu/reg_out[16] ;
 wire \soc/cpu/reg_out[17] ;
 wire \soc/cpu/reg_out[18] ;
 wire \soc/cpu/reg_out[19] ;
 wire \soc/cpu/reg_out[1] ;
 wire \soc/cpu/reg_out[20] ;
 wire \soc/cpu/reg_out[21] ;
 wire \soc/cpu/reg_out[22] ;
 wire \soc/cpu/reg_out[23] ;
 wire \soc/cpu/reg_out[24] ;
 wire \soc/cpu/reg_out[25] ;
 wire \soc/cpu/reg_out[26] ;
 wire \soc/cpu/reg_out[27] ;
 wire \soc/cpu/reg_out[28] ;
 wire \soc/cpu/reg_out[29] ;
 wire \soc/cpu/reg_out[2] ;
 wire \soc/cpu/reg_out[30] ;
 wire \soc/cpu/reg_out[31] ;
 wire \soc/cpu/reg_out[3] ;
 wire \soc/cpu/reg_out[4] ;
 wire \soc/cpu/reg_out[5] ;
 wire \soc/cpu/reg_out[6] ;
 wire \soc/cpu/reg_out[7] ;
 wire \soc/cpu/reg_out[8] ;
 wire \soc/cpu/reg_out[9] ;
 wire \soc/cpu/reg_pc[10] ;
 wire \soc/cpu/reg_pc[11] ;
 wire \soc/cpu/reg_pc[12] ;
 wire \soc/cpu/reg_pc[13] ;
 wire \soc/cpu/reg_pc[14] ;
 wire \soc/cpu/reg_pc[15] ;
 wire \soc/cpu/reg_pc[16] ;
 wire \soc/cpu/reg_pc[17] ;
 wire \soc/cpu/reg_pc[18] ;
 wire \soc/cpu/reg_pc[19] ;
 wire \soc/cpu/reg_pc[1] ;
 wire \soc/cpu/reg_pc[20] ;
 wire \soc/cpu/reg_pc[21] ;
 wire \soc/cpu/reg_pc[22] ;
 wire \soc/cpu/reg_pc[23] ;
 wire \soc/cpu/reg_pc[24] ;
 wire \soc/cpu/reg_pc[25] ;
 wire \soc/cpu/reg_pc[26] ;
 wire \soc/cpu/reg_pc[27] ;
 wire \soc/cpu/reg_pc[28] ;
 wire \soc/cpu/reg_pc[29] ;
 wire \soc/cpu/reg_pc[2] ;
 wire \soc/cpu/reg_pc[30] ;
 wire \soc/cpu/reg_pc[31] ;
 wire \soc/cpu/reg_pc[3] ;
 wire \soc/cpu/reg_pc[4] ;
 wire \soc/cpu/reg_pc[5] ;
 wire \soc/cpu/reg_pc[6] ;
 wire \soc/cpu/reg_pc[7] ;
 wire \soc/cpu/reg_pc[8] ;
 wire \soc/cpu/reg_pc[9] ;
 wire \soc/cpu/reg_sh[0] ;
 wire \soc/cpu/reg_sh[1] ;
 wire \soc/cpu/reg_sh[2] ;
 wire \soc/cpu/reg_sh[3] ;
 wire \soc/cpu/reg_sh[4] ;
 wire \soc/cpu/timer[0] ;
 wire \soc/cpu/timer[10] ;
 wire \soc/cpu/timer[11] ;
 wire \soc/cpu/timer[12] ;
 wire \soc/cpu/timer[13] ;
 wire \soc/cpu/timer[14] ;
 wire \soc/cpu/timer[15] ;
 wire \soc/cpu/timer[16] ;
 wire \soc/cpu/timer[17] ;
 wire \soc/cpu/timer[18] ;
 wire \soc/cpu/timer[19] ;
 wire \soc/cpu/timer[1] ;
 wire \soc/cpu/timer[20] ;
 wire \soc/cpu/timer[21] ;
 wire \soc/cpu/timer[22] ;
 wire \soc/cpu/timer[23] ;
 wire \soc/cpu/timer[24] ;
 wire \soc/cpu/timer[25] ;
 wire \soc/cpu/timer[26] ;
 wire \soc/cpu/timer[27] ;
 wire \soc/cpu/timer[28] ;
 wire \soc/cpu/timer[29] ;
 wire \soc/cpu/timer[2] ;
 wire \soc/cpu/timer[30] ;
 wire \soc/cpu/timer[31] ;
 wire \soc/cpu/timer[3] ;
 wire \soc/cpu/timer[4] ;
 wire \soc/cpu/timer[5] ;
 wire \soc/cpu/timer[6] ;
 wire \soc/cpu/timer[7] ;
 wire \soc/cpu/timer[8] ;
 wire \soc/cpu/timer[9] ;
 wire net667;
 wire net657;
 wire net656;
 wire net655;
 wire net654;
 wire net653;
 wire net652;
 wire net651;
 wire net650;
 wire net649;
 wire net648;
 wire net666;
 wire net647;
 wire net646;
 wire net645;
 wire net644;
 wire net643;
 wire net642;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net665;
 wire net637;
 wire net636;
 wire net635;
 wire net634;
 wire net633;
 wire net632;
 wire net664;
 wire net663;
 wire net662;
 wire net661;
 wire net660;
 wire net659;
 wire net658;
 wire net631;
 wire \soc/cpu/trap ;
 wire \soc/cpu/cpuregs/_0000_ ;
 wire \soc/cpu/cpuregs/_0001_ ;
 wire \soc/cpu/cpuregs/_0002_ ;
 wire \soc/cpu/cpuregs/_0003_ ;
 wire \soc/cpu/cpuregs/_0004_ ;
 wire \soc/cpu/cpuregs/_0005_ ;
 wire \soc/cpu/cpuregs/_0006_ ;
 wire \soc/cpu/cpuregs/_0007_ ;
 wire \soc/cpu/cpuregs/_0008_ ;
 wire \soc/cpu/cpuregs/_0009_ ;
 wire \soc/cpu/cpuregs/_0010_ ;
 wire \soc/cpu/cpuregs/_0011_ ;
 wire \soc/cpu/cpuregs/_0012_ ;
 wire \soc/cpu/cpuregs/_0013_ ;
 wire \soc/cpu/cpuregs/_0014_ ;
 wire \soc/cpu/cpuregs/_0015_ ;
 wire \soc/cpu/cpuregs/_0016_ ;
 wire \soc/cpu/cpuregs/_0017_ ;
 wire \soc/cpu/cpuregs/_0018_ ;
 wire \soc/cpu/cpuregs/_0019_ ;
 wire \soc/cpu/cpuregs/_0020_ ;
 wire \soc/cpu/cpuregs/_0021_ ;
 wire \soc/cpu/cpuregs/_0022_ ;
 wire \soc/cpu/cpuregs/_0023_ ;
 wire \soc/cpu/cpuregs/_0024_ ;
 wire \soc/cpu/cpuregs/_0025_ ;
 wire \soc/cpu/cpuregs/_0026_ ;
 wire \soc/cpu/cpuregs/_0027_ ;
 wire \soc/cpu/cpuregs/_0028_ ;
 wire \soc/cpu/cpuregs/_0029_ ;
 wire \soc/cpu/cpuregs/_0030_ ;
 wire \soc/cpu/cpuregs/_0031_ ;
 wire \soc/cpu/cpuregs/_0032_ ;
 wire \soc/cpu/cpuregs/_0033_ ;
 wire \soc/cpu/cpuregs/_0034_ ;
 wire \soc/cpu/cpuregs/_0035_ ;
 wire \soc/cpu/cpuregs/_0036_ ;
 wire \soc/cpu/cpuregs/_0037_ ;
 wire \soc/cpu/cpuregs/_0038_ ;
 wire \soc/cpu/cpuregs/_0039_ ;
 wire \soc/cpu/cpuregs/_0040_ ;
 wire \soc/cpu/cpuregs/_0041_ ;
 wire \soc/cpu/cpuregs/_0042_ ;
 wire \soc/cpu/cpuregs/_0043_ ;
 wire \soc/cpu/cpuregs/_0044_ ;
 wire \soc/cpu/cpuregs/_0045_ ;
 wire \soc/cpu/cpuregs/_0046_ ;
 wire \soc/cpu/cpuregs/_0047_ ;
 wire \soc/cpu/cpuregs/_0048_ ;
 wire \soc/cpu/cpuregs/_0049_ ;
 wire \soc/cpu/cpuregs/_0050_ ;
 wire \soc/cpu/cpuregs/_0051_ ;
 wire \soc/cpu/cpuregs/_0052_ ;
 wire \soc/cpu/cpuregs/_0053_ ;
 wire \soc/cpu/cpuregs/_0054_ ;
 wire \soc/cpu/cpuregs/_0055_ ;
 wire \soc/cpu/cpuregs/_0056_ ;
 wire \soc/cpu/cpuregs/_0057_ ;
 wire \soc/cpu/cpuregs/_0058_ ;
 wire \soc/cpu/cpuregs/_0059_ ;
 wire \soc/cpu/cpuregs/_0060_ ;
 wire \soc/cpu/cpuregs/_0061_ ;
 wire \soc/cpu/cpuregs/_0062_ ;
 wire \soc/cpu/cpuregs/_0063_ ;
 wire \soc/cpu/cpuregs/_0064_ ;
 wire \soc/cpu/cpuregs/_0065_ ;
 wire \soc/cpu/cpuregs/_0066_ ;
 wire \soc/cpu/cpuregs/_0067_ ;
 wire \soc/cpu/cpuregs/_0068_ ;
 wire \soc/cpu/cpuregs/_0069_ ;
 wire \soc/cpu/cpuregs/_0070_ ;
 wire \soc/cpu/cpuregs/_0071_ ;
 wire \soc/cpu/cpuregs/_0072_ ;
 wire \soc/cpu/cpuregs/_0073_ ;
 wire \soc/cpu/cpuregs/_0074_ ;
 wire \soc/cpu/cpuregs/_0075_ ;
 wire \soc/cpu/cpuregs/_0076_ ;
 wire \soc/cpu/cpuregs/_0077_ ;
 wire \soc/cpu/cpuregs/_0078_ ;
 wire \soc/cpu/cpuregs/_0079_ ;
 wire \soc/cpu/cpuregs/_0080_ ;
 wire \soc/cpu/cpuregs/_0081_ ;
 wire \soc/cpu/cpuregs/_0082_ ;
 wire \soc/cpu/cpuregs/_0083_ ;
 wire \soc/cpu/cpuregs/_0084_ ;
 wire \soc/cpu/cpuregs/_0085_ ;
 wire \soc/cpu/cpuregs/_0086_ ;
 wire \soc/cpu/cpuregs/_0087_ ;
 wire \soc/cpu/cpuregs/_0088_ ;
 wire \soc/cpu/cpuregs/_0089_ ;
 wire \soc/cpu/cpuregs/_0090_ ;
 wire \soc/cpu/cpuregs/_0091_ ;
 wire \soc/cpu/cpuregs/_0092_ ;
 wire \soc/cpu/cpuregs/_0093_ ;
 wire \soc/cpu/cpuregs/_0094_ ;
 wire \soc/cpu/cpuregs/_0095_ ;
 wire \soc/cpu/cpuregs/_0096_ ;
 wire \soc/cpu/cpuregs/_0097_ ;
 wire \soc/cpu/cpuregs/_0098_ ;
 wire \soc/cpu/cpuregs/_0099_ ;
 wire \soc/cpu/cpuregs/_0100_ ;
 wire \soc/cpu/cpuregs/_0101_ ;
 wire \soc/cpu/cpuregs/_0102_ ;
 wire \soc/cpu/cpuregs/_0103_ ;
 wire \soc/cpu/cpuregs/_0104_ ;
 wire \soc/cpu/cpuregs/_0105_ ;
 wire \soc/cpu/cpuregs/_0106_ ;
 wire \soc/cpu/cpuregs/_0107_ ;
 wire \soc/cpu/cpuregs/_0108_ ;
 wire \soc/cpu/cpuregs/_0109_ ;
 wire \soc/cpu/cpuregs/_0110_ ;
 wire \soc/cpu/cpuregs/_0111_ ;
 wire \soc/cpu/cpuregs/_0112_ ;
 wire \soc/cpu/cpuregs/_0113_ ;
 wire \soc/cpu/cpuregs/_0114_ ;
 wire \soc/cpu/cpuregs/_0115_ ;
 wire \soc/cpu/cpuregs/_0116_ ;
 wire \soc/cpu/cpuregs/_0117_ ;
 wire \soc/cpu/cpuregs/_0118_ ;
 wire \soc/cpu/cpuregs/_0119_ ;
 wire \soc/cpu/cpuregs/_0120_ ;
 wire \soc/cpu/cpuregs/_0121_ ;
 wire \soc/cpu/cpuregs/_0122_ ;
 wire \soc/cpu/cpuregs/_0123_ ;
 wire \soc/cpu/cpuregs/_0124_ ;
 wire \soc/cpu/cpuregs/_0125_ ;
 wire \soc/cpu/cpuregs/_0126_ ;
 wire \soc/cpu/cpuregs/_0127_ ;
 wire \soc/cpu/cpuregs/_0128_ ;
 wire \soc/cpu/cpuregs/_0129_ ;
 wire \soc/cpu/cpuregs/_0130_ ;
 wire \soc/cpu/cpuregs/_0131_ ;
 wire \soc/cpu/cpuregs/_0132_ ;
 wire \soc/cpu/cpuregs/_0133_ ;
 wire \soc/cpu/cpuregs/_0134_ ;
 wire \soc/cpu/cpuregs/_0135_ ;
 wire \soc/cpu/cpuregs/_0136_ ;
 wire \soc/cpu/cpuregs/_0137_ ;
 wire \soc/cpu/cpuregs/_0138_ ;
 wire \soc/cpu/cpuregs/_0139_ ;
 wire \soc/cpu/cpuregs/_0140_ ;
 wire \soc/cpu/cpuregs/_0141_ ;
 wire \soc/cpu/cpuregs/_0142_ ;
 wire \soc/cpu/cpuregs/_0143_ ;
 wire \soc/cpu/cpuregs/_0144_ ;
 wire \soc/cpu/cpuregs/_0145_ ;
 wire \soc/cpu/cpuregs/_0146_ ;
 wire \soc/cpu/cpuregs/_0147_ ;
 wire \soc/cpu/cpuregs/_0148_ ;
 wire \soc/cpu/cpuregs/_0149_ ;
 wire \soc/cpu/cpuregs/_0150_ ;
 wire \soc/cpu/cpuregs/_0151_ ;
 wire \soc/cpu/cpuregs/_0152_ ;
 wire \soc/cpu/cpuregs/_0153_ ;
 wire \soc/cpu/cpuregs/_0154_ ;
 wire \soc/cpu/cpuregs/_0155_ ;
 wire \soc/cpu/cpuregs/_0156_ ;
 wire \soc/cpu/cpuregs/_0157_ ;
 wire \soc/cpu/cpuregs/_0158_ ;
 wire \soc/cpu/cpuregs/_0159_ ;
 wire \soc/cpu/cpuregs/_0160_ ;
 wire \soc/cpu/cpuregs/_0161_ ;
 wire \soc/cpu/cpuregs/_0162_ ;
 wire \soc/cpu/cpuregs/_0163_ ;
 wire \soc/cpu/cpuregs/_0164_ ;
 wire \soc/cpu/cpuregs/_0165_ ;
 wire \soc/cpu/cpuregs/_0166_ ;
 wire \soc/cpu/cpuregs/_0167_ ;
 wire \soc/cpu/cpuregs/_0168_ ;
 wire \soc/cpu/cpuregs/_0169_ ;
 wire \soc/cpu/cpuregs/_0170_ ;
 wire \soc/cpu/cpuregs/_0171_ ;
 wire \soc/cpu/cpuregs/_0172_ ;
 wire \soc/cpu/cpuregs/_0173_ ;
 wire \soc/cpu/cpuregs/_0174_ ;
 wire \soc/cpu/cpuregs/_0175_ ;
 wire \soc/cpu/cpuregs/_0176_ ;
 wire \soc/cpu/cpuregs/_0177_ ;
 wire \soc/cpu/cpuregs/_0178_ ;
 wire \soc/cpu/cpuregs/_0179_ ;
 wire \soc/cpu/cpuregs/_0180_ ;
 wire \soc/cpu/cpuregs/_0181_ ;
 wire \soc/cpu/cpuregs/_0182_ ;
 wire \soc/cpu/cpuregs/_0183_ ;
 wire \soc/cpu/cpuregs/_0184_ ;
 wire \soc/cpu/cpuregs/_0185_ ;
 wire \soc/cpu/cpuregs/_0186_ ;
 wire \soc/cpu/cpuregs/_0187_ ;
 wire \soc/cpu/cpuregs/_0188_ ;
 wire \soc/cpu/cpuregs/_0189_ ;
 wire \soc/cpu/cpuregs/_0190_ ;
 wire \soc/cpu/cpuregs/_0191_ ;
 wire \soc/cpu/cpuregs/_0192_ ;
 wire \soc/cpu/cpuregs/_0193_ ;
 wire \soc/cpu/cpuregs/_0194_ ;
 wire \soc/cpu/cpuregs/_0195_ ;
 wire \soc/cpu/cpuregs/_0196_ ;
 wire \soc/cpu/cpuregs/_0197_ ;
 wire \soc/cpu/cpuregs/_0198_ ;
 wire \soc/cpu/cpuregs/_0199_ ;
 wire \soc/cpu/cpuregs/_0200_ ;
 wire \soc/cpu/cpuregs/_0201_ ;
 wire \soc/cpu/cpuregs/_0202_ ;
 wire \soc/cpu/cpuregs/_0203_ ;
 wire \soc/cpu/cpuregs/_0204_ ;
 wire \soc/cpu/cpuregs/_0205_ ;
 wire \soc/cpu/cpuregs/_0206_ ;
 wire \soc/cpu/cpuregs/_0207_ ;
 wire \soc/cpu/cpuregs/_0208_ ;
 wire \soc/cpu/cpuregs/_0209_ ;
 wire \soc/cpu/cpuregs/_0210_ ;
 wire \soc/cpu/cpuregs/_0211_ ;
 wire \soc/cpu/cpuregs/_0212_ ;
 wire \soc/cpu/cpuregs/_0213_ ;
 wire \soc/cpu/cpuregs/_0214_ ;
 wire \soc/cpu/cpuregs/_0215_ ;
 wire \soc/cpu/cpuregs/_0216_ ;
 wire \soc/cpu/cpuregs/_0217_ ;
 wire \soc/cpu/cpuregs/_0218_ ;
 wire \soc/cpu/cpuregs/_0219_ ;
 wire \soc/cpu/cpuregs/_0220_ ;
 wire \soc/cpu/cpuregs/_0221_ ;
 wire \soc/cpu/cpuregs/_0222_ ;
 wire \soc/cpu/cpuregs/_0223_ ;
 wire \soc/cpu/cpuregs/_0224_ ;
 wire \soc/cpu/cpuregs/_0225_ ;
 wire \soc/cpu/cpuregs/_0226_ ;
 wire \soc/cpu/cpuregs/_0227_ ;
 wire \soc/cpu/cpuregs/_0228_ ;
 wire \soc/cpu/cpuregs/_0229_ ;
 wire \soc/cpu/cpuregs/_0230_ ;
 wire \soc/cpu/cpuregs/_0231_ ;
 wire \soc/cpu/cpuregs/_0232_ ;
 wire \soc/cpu/cpuregs/_0233_ ;
 wire \soc/cpu/cpuregs/_0234_ ;
 wire \soc/cpu/cpuregs/_0235_ ;
 wire \soc/cpu/cpuregs/_0236_ ;
 wire \soc/cpu/cpuregs/_0237_ ;
 wire \soc/cpu/cpuregs/_0238_ ;
 wire \soc/cpu/cpuregs/_0239_ ;
 wire \soc/cpu/cpuregs/_0240_ ;
 wire \soc/cpu/cpuregs/_0241_ ;
 wire \soc/cpu/cpuregs/_0242_ ;
 wire \soc/cpu/cpuregs/_0243_ ;
 wire \soc/cpu/cpuregs/_0244_ ;
 wire \soc/cpu/cpuregs/_0245_ ;
 wire \soc/cpu/cpuregs/_0246_ ;
 wire \soc/cpu/cpuregs/_0247_ ;
 wire \soc/cpu/cpuregs/_0248_ ;
 wire \soc/cpu/cpuregs/_0249_ ;
 wire \soc/cpu/cpuregs/_0250_ ;
 wire \soc/cpu/cpuregs/_0251_ ;
 wire \soc/cpu/cpuregs/_0252_ ;
 wire \soc/cpu/cpuregs/_0253_ ;
 wire \soc/cpu/cpuregs/_0254_ ;
 wire \soc/cpu/cpuregs/_0255_ ;
 wire \soc/cpu/cpuregs/_0256_ ;
 wire \soc/cpu/cpuregs/_0257_ ;
 wire \soc/cpu/cpuregs/_0258_ ;
 wire \soc/cpu/cpuregs/_0259_ ;
 wire \soc/cpu/cpuregs/_0260_ ;
 wire \soc/cpu/cpuregs/_0261_ ;
 wire \soc/cpu/cpuregs/_0262_ ;
 wire \soc/cpu/cpuregs/_0263_ ;
 wire \soc/cpu/cpuregs/_0264_ ;
 wire \soc/cpu/cpuregs/_0265_ ;
 wire \soc/cpu/cpuregs/_0266_ ;
 wire \soc/cpu/cpuregs/_0267_ ;
 wire \soc/cpu/cpuregs/_0268_ ;
 wire \soc/cpu/cpuregs/_0269_ ;
 wire \soc/cpu/cpuregs/_0270_ ;
 wire \soc/cpu/cpuregs/_0271_ ;
 wire \soc/cpu/cpuregs/_0272_ ;
 wire \soc/cpu/cpuregs/_0273_ ;
 wire \soc/cpu/cpuregs/_0274_ ;
 wire \soc/cpu/cpuregs/_0275_ ;
 wire \soc/cpu/cpuregs/_0276_ ;
 wire \soc/cpu/cpuregs/_0277_ ;
 wire \soc/cpu/cpuregs/_0278_ ;
 wire \soc/cpu/cpuregs/_0279_ ;
 wire \soc/cpu/cpuregs/_0280_ ;
 wire \soc/cpu/cpuregs/_0281_ ;
 wire \soc/cpu/cpuregs/_0282_ ;
 wire \soc/cpu/cpuregs/_0283_ ;
 wire \soc/cpu/cpuregs/_0284_ ;
 wire \soc/cpu/cpuregs/_0285_ ;
 wire \soc/cpu/cpuregs/_0286_ ;
 wire \soc/cpu/cpuregs/_0287_ ;
 wire \soc/cpu/cpuregs/_0288_ ;
 wire \soc/cpu/cpuregs/_0289_ ;
 wire \soc/cpu/cpuregs/_0290_ ;
 wire \soc/cpu/cpuregs/_0291_ ;
 wire \soc/cpu/cpuregs/_0292_ ;
 wire \soc/cpu/cpuregs/_0293_ ;
 wire \soc/cpu/cpuregs/_0294_ ;
 wire \soc/cpu/cpuregs/_0295_ ;
 wire \soc/cpu/cpuregs/_0296_ ;
 wire \soc/cpu/cpuregs/_0297_ ;
 wire \soc/cpu/cpuregs/_0298_ ;
 wire \soc/cpu/cpuregs/_0299_ ;
 wire \soc/cpu/cpuregs/_0300_ ;
 wire \soc/cpu/cpuregs/_0301_ ;
 wire \soc/cpu/cpuregs/_0302_ ;
 wire \soc/cpu/cpuregs/_0303_ ;
 wire \soc/cpu/cpuregs/_0304_ ;
 wire \soc/cpu/cpuregs/_0305_ ;
 wire \soc/cpu/cpuregs/_0306_ ;
 wire \soc/cpu/cpuregs/_0307_ ;
 wire \soc/cpu/cpuregs/_0308_ ;
 wire \soc/cpu/cpuregs/_0309_ ;
 wire \soc/cpu/cpuregs/_0310_ ;
 wire \soc/cpu/cpuregs/_0311_ ;
 wire \soc/cpu/cpuregs/_0312_ ;
 wire \soc/cpu/cpuregs/_0313_ ;
 wire \soc/cpu/cpuregs/_0314_ ;
 wire \soc/cpu/cpuregs/_0315_ ;
 wire \soc/cpu/cpuregs/_0316_ ;
 wire \soc/cpu/cpuregs/_0317_ ;
 wire \soc/cpu/cpuregs/_0318_ ;
 wire \soc/cpu/cpuregs/_0319_ ;
 wire \soc/cpu/cpuregs/_0320_ ;
 wire \soc/cpu/cpuregs/_0321_ ;
 wire \soc/cpu/cpuregs/_0322_ ;
 wire \soc/cpu/cpuregs/_0323_ ;
 wire \soc/cpu/cpuregs/_0324_ ;
 wire \soc/cpu/cpuregs/_0325_ ;
 wire \soc/cpu/cpuregs/_0326_ ;
 wire \soc/cpu/cpuregs/_0327_ ;
 wire \soc/cpu/cpuregs/_0328_ ;
 wire \soc/cpu/cpuregs/_0329_ ;
 wire \soc/cpu/cpuregs/_0330_ ;
 wire \soc/cpu/cpuregs/_0331_ ;
 wire \soc/cpu/cpuregs/_0332_ ;
 wire \soc/cpu/cpuregs/_0333_ ;
 wire \soc/cpu/cpuregs/_0334_ ;
 wire \soc/cpu/cpuregs/_0335_ ;
 wire \soc/cpu/cpuregs/_0336_ ;
 wire \soc/cpu/cpuregs/_0337_ ;
 wire \soc/cpu/cpuregs/_0338_ ;
 wire \soc/cpu/cpuregs/_0339_ ;
 wire \soc/cpu/cpuregs/_0340_ ;
 wire \soc/cpu/cpuregs/_0341_ ;
 wire \soc/cpu/cpuregs/_0342_ ;
 wire \soc/cpu/cpuregs/_0343_ ;
 wire \soc/cpu/cpuregs/_0344_ ;
 wire \soc/cpu/cpuregs/_0345_ ;
 wire \soc/cpu/cpuregs/_0346_ ;
 wire \soc/cpu/cpuregs/_0347_ ;
 wire \soc/cpu/cpuregs/_0348_ ;
 wire \soc/cpu/cpuregs/_0349_ ;
 wire \soc/cpu/cpuregs/_0350_ ;
 wire \soc/cpu/cpuregs/_0351_ ;
 wire \soc/cpu/cpuregs/_0352_ ;
 wire \soc/cpu/cpuregs/_0353_ ;
 wire \soc/cpu/cpuregs/_0354_ ;
 wire \soc/cpu/cpuregs/_0355_ ;
 wire \soc/cpu/cpuregs/_0356_ ;
 wire \soc/cpu/cpuregs/_0357_ ;
 wire \soc/cpu/cpuregs/_0358_ ;
 wire \soc/cpu/cpuregs/_0359_ ;
 wire \soc/cpu/cpuregs/_0360_ ;
 wire \soc/cpu/cpuregs/_0361_ ;
 wire \soc/cpu/cpuregs/_0362_ ;
 wire \soc/cpu/cpuregs/_0363_ ;
 wire \soc/cpu/cpuregs/_0364_ ;
 wire \soc/cpu/cpuregs/_0365_ ;
 wire \soc/cpu/cpuregs/_0366_ ;
 wire \soc/cpu/cpuregs/_0367_ ;
 wire \soc/cpu/cpuregs/_0368_ ;
 wire \soc/cpu/cpuregs/_0369_ ;
 wire \soc/cpu/cpuregs/_0370_ ;
 wire \soc/cpu/cpuregs/_0371_ ;
 wire \soc/cpu/cpuregs/_0372_ ;
 wire \soc/cpu/cpuregs/_0373_ ;
 wire \soc/cpu/cpuregs/_0374_ ;
 wire \soc/cpu/cpuregs/_0375_ ;
 wire \soc/cpu/cpuregs/_0376_ ;
 wire \soc/cpu/cpuregs/_0377_ ;
 wire \soc/cpu/cpuregs/_0378_ ;
 wire \soc/cpu/cpuregs/_0379_ ;
 wire \soc/cpu/cpuregs/_0380_ ;
 wire \soc/cpu/cpuregs/_0381_ ;
 wire \soc/cpu/cpuregs/_0382_ ;
 wire \soc/cpu/cpuregs/_0383_ ;
 wire \soc/cpu/cpuregs/_0384_ ;
 wire \soc/cpu/cpuregs/_0385_ ;
 wire \soc/cpu/cpuregs/_0386_ ;
 wire \soc/cpu/cpuregs/_0387_ ;
 wire \soc/cpu/cpuregs/_0388_ ;
 wire \soc/cpu/cpuregs/_0389_ ;
 wire \soc/cpu/cpuregs/_0390_ ;
 wire \soc/cpu/cpuregs/_0391_ ;
 wire \soc/cpu/cpuregs/_0392_ ;
 wire \soc/cpu/cpuregs/_0393_ ;
 wire \soc/cpu/cpuregs/_0394_ ;
 wire \soc/cpu/cpuregs/_0395_ ;
 wire \soc/cpu/cpuregs/_0396_ ;
 wire \soc/cpu/cpuregs/_0397_ ;
 wire \soc/cpu/cpuregs/_0398_ ;
 wire \soc/cpu/cpuregs/_0399_ ;
 wire \soc/cpu/cpuregs/_0400_ ;
 wire \soc/cpu/cpuregs/_0401_ ;
 wire \soc/cpu/cpuregs/_0402_ ;
 wire \soc/cpu/cpuregs/_0403_ ;
 wire \soc/cpu/cpuregs/_0404_ ;
 wire \soc/cpu/cpuregs/_0405_ ;
 wire \soc/cpu/cpuregs/_0406_ ;
 wire \soc/cpu/cpuregs/_0407_ ;
 wire \soc/cpu/cpuregs/_0408_ ;
 wire \soc/cpu/cpuregs/_0409_ ;
 wire \soc/cpu/cpuregs/_0410_ ;
 wire \soc/cpu/cpuregs/_0411_ ;
 wire \soc/cpu/cpuregs/_0412_ ;
 wire \soc/cpu/cpuregs/_0413_ ;
 wire \soc/cpu/cpuregs/_0414_ ;
 wire \soc/cpu/cpuregs/_0415_ ;
 wire \soc/cpu/cpuregs/_0416_ ;
 wire \soc/cpu/cpuregs/_0417_ ;
 wire \soc/cpu/cpuregs/_0418_ ;
 wire \soc/cpu/cpuregs/_0419_ ;
 wire \soc/cpu/cpuregs/_0420_ ;
 wire \soc/cpu/cpuregs/_0421_ ;
 wire \soc/cpu/cpuregs/_0422_ ;
 wire \soc/cpu/cpuregs/_0423_ ;
 wire \soc/cpu/cpuregs/_0424_ ;
 wire \soc/cpu/cpuregs/_0425_ ;
 wire \soc/cpu/cpuregs/_0426_ ;
 wire \soc/cpu/cpuregs/_0427_ ;
 wire \soc/cpu/cpuregs/_0428_ ;
 wire \soc/cpu/cpuregs/_0429_ ;
 wire \soc/cpu/cpuregs/_0430_ ;
 wire \soc/cpu/cpuregs/_0431_ ;
 wire \soc/cpu/cpuregs/_0432_ ;
 wire \soc/cpu/cpuregs/_0433_ ;
 wire \soc/cpu/cpuregs/_0434_ ;
 wire \soc/cpu/cpuregs/_0435_ ;
 wire \soc/cpu/cpuregs/_0436_ ;
 wire \soc/cpu/cpuregs/_0437_ ;
 wire \soc/cpu/cpuregs/_0438_ ;
 wire \soc/cpu/cpuregs/_0439_ ;
 wire \soc/cpu/cpuregs/_0440_ ;
 wire \soc/cpu/cpuregs/_0441_ ;
 wire \soc/cpu/cpuregs/_0442_ ;
 wire \soc/cpu/cpuregs/_0443_ ;
 wire \soc/cpu/cpuregs/_0444_ ;
 wire \soc/cpu/cpuregs/_0445_ ;
 wire \soc/cpu/cpuregs/_0446_ ;
 wire \soc/cpu/cpuregs/_0447_ ;
 wire \soc/cpu/cpuregs/_0448_ ;
 wire \soc/cpu/cpuregs/_0449_ ;
 wire \soc/cpu/cpuregs/_0450_ ;
 wire \soc/cpu/cpuregs/_0451_ ;
 wire \soc/cpu/cpuregs/_0452_ ;
 wire \soc/cpu/cpuregs/_0453_ ;
 wire \soc/cpu/cpuregs/_0454_ ;
 wire \soc/cpu/cpuregs/_0455_ ;
 wire \soc/cpu/cpuregs/_0456_ ;
 wire \soc/cpu/cpuregs/_0457_ ;
 wire \soc/cpu/cpuregs/_0458_ ;
 wire \soc/cpu/cpuregs/_0459_ ;
 wire \soc/cpu/cpuregs/_0460_ ;
 wire \soc/cpu/cpuregs/_0461_ ;
 wire \soc/cpu/cpuregs/_0462_ ;
 wire \soc/cpu/cpuregs/_0463_ ;
 wire \soc/cpu/cpuregs/_0464_ ;
 wire \soc/cpu/cpuregs/_0465_ ;
 wire \soc/cpu/cpuregs/_0466_ ;
 wire \soc/cpu/cpuregs/_0467_ ;
 wire \soc/cpu/cpuregs/_0468_ ;
 wire \soc/cpu/cpuregs/_0469_ ;
 wire \soc/cpu/cpuregs/_0470_ ;
 wire \soc/cpu/cpuregs/_0471_ ;
 wire \soc/cpu/cpuregs/_0472_ ;
 wire \soc/cpu/cpuregs/_0473_ ;
 wire \soc/cpu/cpuregs/_0474_ ;
 wire \soc/cpu/cpuregs/_0475_ ;
 wire \soc/cpu/cpuregs/_0476_ ;
 wire \soc/cpu/cpuregs/_0477_ ;
 wire \soc/cpu/cpuregs/_0478_ ;
 wire \soc/cpu/cpuregs/_0479_ ;
 wire \soc/cpu/cpuregs/_0480_ ;
 wire \soc/cpu/cpuregs/_0481_ ;
 wire \soc/cpu/cpuregs/_0482_ ;
 wire \soc/cpu/cpuregs/_0483_ ;
 wire \soc/cpu/cpuregs/_0484_ ;
 wire \soc/cpu/cpuregs/_0485_ ;
 wire \soc/cpu/cpuregs/_0486_ ;
 wire \soc/cpu/cpuregs/_0487_ ;
 wire \soc/cpu/cpuregs/_0488_ ;
 wire \soc/cpu/cpuregs/_0489_ ;
 wire \soc/cpu/cpuregs/_0490_ ;
 wire \soc/cpu/cpuregs/_0491_ ;
 wire \soc/cpu/cpuregs/_0492_ ;
 wire \soc/cpu/cpuregs/_0493_ ;
 wire \soc/cpu/cpuregs/_0494_ ;
 wire \soc/cpu/cpuregs/_0495_ ;
 wire \soc/cpu/cpuregs/_0496_ ;
 wire \soc/cpu/cpuregs/_0497_ ;
 wire \soc/cpu/cpuregs/_0498_ ;
 wire \soc/cpu/cpuregs/_0499_ ;
 wire \soc/cpu/cpuregs/_0500_ ;
 wire \soc/cpu/cpuregs/_0501_ ;
 wire \soc/cpu/cpuregs/_0502_ ;
 wire \soc/cpu/cpuregs/_0503_ ;
 wire \soc/cpu/cpuregs/_0504_ ;
 wire \soc/cpu/cpuregs/_0505_ ;
 wire \soc/cpu/cpuregs/_0506_ ;
 wire \soc/cpu/cpuregs/_0507_ ;
 wire \soc/cpu/cpuregs/_0508_ ;
 wire \soc/cpu/cpuregs/_0509_ ;
 wire \soc/cpu/cpuregs/_0510_ ;
 wire \soc/cpu/cpuregs/_0511_ ;
 wire \soc/cpu/cpuregs/_0512_ ;
 wire \soc/cpu/cpuregs/_0513_ ;
 wire \soc/cpu/cpuregs/_0514_ ;
 wire \soc/cpu/cpuregs/_0515_ ;
 wire \soc/cpu/cpuregs/_0516_ ;
 wire \soc/cpu/cpuregs/_0517_ ;
 wire \soc/cpu/cpuregs/_0518_ ;
 wire \soc/cpu/cpuregs/_0519_ ;
 wire \soc/cpu/cpuregs/_0520_ ;
 wire \soc/cpu/cpuregs/_0521_ ;
 wire \soc/cpu/cpuregs/_0522_ ;
 wire \soc/cpu/cpuregs/_0523_ ;
 wire \soc/cpu/cpuregs/_0524_ ;
 wire \soc/cpu/cpuregs/_0525_ ;
 wire \soc/cpu/cpuregs/_0526_ ;
 wire \soc/cpu/cpuregs/_0527_ ;
 wire \soc/cpu/cpuregs/_0528_ ;
 wire \soc/cpu/cpuregs/_0529_ ;
 wire \soc/cpu/cpuregs/_0530_ ;
 wire \soc/cpu/cpuregs/_0531_ ;
 wire \soc/cpu/cpuregs/_0532_ ;
 wire \soc/cpu/cpuregs/_0533_ ;
 wire \soc/cpu/cpuregs/_0534_ ;
 wire \soc/cpu/cpuregs/_0535_ ;
 wire \soc/cpu/cpuregs/_0536_ ;
 wire \soc/cpu/cpuregs/_0537_ ;
 wire \soc/cpu/cpuregs/_0538_ ;
 wire \soc/cpu/cpuregs/_0539_ ;
 wire \soc/cpu/cpuregs/_0540_ ;
 wire \soc/cpu/cpuregs/_0541_ ;
 wire \soc/cpu/cpuregs/_0542_ ;
 wire \soc/cpu/cpuregs/_0543_ ;
 wire \soc/cpu/cpuregs/_0544_ ;
 wire \soc/cpu/cpuregs/_0545_ ;
 wire \soc/cpu/cpuregs/_0546_ ;
 wire \soc/cpu/cpuregs/_0547_ ;
 wire \soc/cpu/cpuregs/_0548_ ;
 wire \soc/cpu/cpuregs/_0549_ ;
 wire \soc/cpu/cpuregs/_0550_ ;
 wire \soc/cpu/cpuregs/_0551_ ;
 wire \soc/cpu/cpuregs/_0552_ ;
 wire \soc/cpu/cpuregs/_0553_ ;
 wire \soc/cpu/cpuregs/_0554_ ;
 wire \soc/cpu/cpuregs/_0555_ ;
 wire \soc/cpu/cpuregs/_0556_ ;
 wire \soc/cpu/cpuregs/_0557_ ;
 wire \soc/cpu/cpuregs/_0558_ ;
 wire \soc/cpu/cpuregs/_0559_ ;
 wire \soc/cpu/cpuregs/_0560_ ;
 wire \soc/cpu/cpuregs/_0561_ ;
 wire \soc/cpu/cpuregs/_0562_ ;
 wire \soc/cpu/cpuregs/_0563_ ;
 wire \soc/cpu/cpuregs/_0564_ ;
 wire \soc/cpu/cpuregs/_0565_ ;
 wire \soc/cpu/cpuregs/_0566_ ;
 wire \soc/cpu/cpuregs/_0567_ ;
 wire \soc/cpu/cpuregs/_0568_ ;
 wire \soc/cpu/cpuregs/_0569_ ;
 wire \soc/cpu/cpuregs/_0570_ ;
 wire \soc/cpu/cpuregs/_0571_ ;
 wire \soc/cpu/cpuregs/_0572_ ;
 wire \soc/cpu/cpuregs/_0573_ ;
 wire \soc/cpu/cpuregs/_0574_ ;
 wire \soc/cpu/cpuregs/_0575_ ;
 wire \soc/cpu/cpuregs/_0576_ ;
 wire \soc/cpu/cpuregs/_0577_ ;
 wire \soc/cpu/cpuregs/_0578_ ;
 wire \soc/cpu/cpuregs/_0579_ ;
 wire \soc/cpu/cpuregs/_0580_ ;
 wire \soc/cpu/cpuregs/_0581_ ;
 wire \soc/cpu/cpuregs/_0582_ ;
 wire \soc/cpu/cpuregs/_0583_ ;
 wire \soc/cpu/cpuregs/_0584_ ;
 wire \soc/cpu/cpuregs/_0585_ ;
 wire \soc/cpu/cpuregs/_0586_ ;
 wire \soc/cpu/cpuregs/_0587_ ;
 wire \soc/cpu/cpuregs/_0588_ ;
 wire \soc/cpu/cpuregs/_0589_ ;
 wire \soc/cpu/cpuregs/_0590_ ;
 wire \soc/cpu/cpuregs/_0591_ ;
 wire \soc/cpu/cpuregs/_0592_ ;
 wire \soc/cpu/cpuregs/_0593_ ;
 wire \soc/cpu/cpuregs/_0594_ ;
 wire \soc/cpu/cpuregs/_0595_ ;
 wire \soc/cpu/cpuregs/_0596_ ;
 wire \soc/cpu/cpuregs/_0597_ ;
 wire \soc/cpu/cpuregs/_0598_ ;
 wire \soc/cpu/cpuregs/_0599_ ;
 wire \soc/cpu/cpuregs/_0600_ ;
 wire \soc/cpu/cpuregs/_0601_ ;
 wire \soc/cpu/cpuregs/_0602_ ;
 wire \soc/cpu/cpuregs/_0603_ ;
 wire \soc/cpu/cpuregs/_0604_ ;
 wire \soc/cpu/cpuregs/_0605_ ;
 wire \soc/cpu/cpuregs/_0606_ ;
 wire \soc/cpu/cpuregs/_0607_ ;
 wire \soc/cpu/cpuregs/_0608_ ;
 wire \soc/cpu/cpuregs/_0609_ ;
 wire \soc/cpu/cpuregs/_0610_ ;
 wire \soc/cpu/cpuregs/_0611_ ;
 wire \soc/cpu/cpuregs/_0612_ ;
 wire \soc/cpu/cpuregs/_0613_ ;
 wire \soc/cpu/cpuregs/_0614_ ;
 wire \soc/cpu/cpuregs/_0615_ ;
 wire \soc/cpu/cpuregs/_0616_ ;
 wire \soc/cpu/cpuregs/_0617_ ;
 wire \soc/cpu/cpuregs/_0618_ ;
 wire \soc/cpu/cpuregs/_0619_ ;
 wire \soc/cpu/cpuregs/_0620_ ;
 wire \soc/cpu/cpuregs/_0621_ ;
 wire \soc/cpu/cpuregs/_0622_ ;
 wire \soc/cpu/cpuregs/_0623_ ;
 wire \soc/cpu/cpuregs/_0624_ ;
 wire \soc/cpu/cpuregs/_0625_ ;
 wire \soc/cpu/cpuregs/_0626_ ;
 wire \soc/cpu/cpuregs/_0627_ ;
 wire \soc/cpu/cpuregs/_0628_ ;
 wire \soc/cpu/cpuregs/_0629_ ;
 wire \soc/cpu/cpuregs/_0630_ ;
 wire \soc/cpu/cpuregs/_0631_ ;
 wire \soc/cpu/cpuregs/_0632_ ;
 wire \soc/cpu/cpuregs/_0633_ ;
 wire \soc/cpu/cpuregs/_0634_ ;
 wire \soc/cpu/cpuregs/_0635_ ;
 wire \soc/cpu/cpuregs/_0636_ ;
 wire \soc/cpu/cpuregs/_0637_ ;
 wire \soc/cpu/cpuregs/_0638_ ;
 wire \soc/cpu/cpuregs/_0639_ ;
 wire \soc/cpu/cpuregs/_0640_ ;
 wire \soc/cpu/cpuregs/_0641_ ;
 wire \soc/cpu/cpuregs/_0642_ ;
 wire \soc/cpu/cpuregs/_0643_ ;
 wire \soc/cpu/cpuregs/_0644_ ;
 wire \soc/cpu/cpuregs/_0645_ ;
 wire \soc/cpu/cpuregs/_0646_ ;
 wire \soc/cpu/cpuregs/_0647_ ;
 wire \soc/cpu/cpuregs/_0648_ ;
 wire \soc/cpu/cpuregs/_0649_ ;
 wire \soc/cpu/cpuregs/_0650_ ;
 wire \soc/cpu/cpuregs/_0651_ ;
 wire \soc/cpu/cpuregs/_0652_ ;
 wire \soc/cpu/cpuregs/_0653_ ;
 wire \soc/cpu/cpuregs/_0654_ ;
 wire \soc/cpu/cpuregs/_0655_ ;
 wire \soc/cpu/cpuregs/_0656_ ;
 wire \soc/cpu/cpuregs/_0657_ ;
 wire \soc/cpu/cpuregs/_0658_ ;
 wire \soc/cpu/cpuregs/_0659_ ;
 wire \soc/cpu/cpuregs/_0660_ ;
 wire \soc/cpu/cpuregs/_0661_ ;
 wire \soc/cpu/cpuregs/_0662_ ;
 wire \soc/cpu/cpuregs/_0663_ ;
 wire \soc/cpu/cpuregs/_0664_ ;
 wire \soc/cpu/cpuregs/_0665_ ;
 wire \soc/cpu/cpuregs/_0666_ ;
 wire \soc/cpu/cpuregs/_0667_ ;
 wire \soc/cpu/cpuregs/_0668_ ;
 wire \soc/cpu/cpuregs/_0669_ ;
 wire \soc/cpu/cpuregs/_0670_ ;
 wire \soc/cpu/cpuregs/_0671_ ;
 wire \soc/cpu/cpuregs/_0672_ ;
 wire \soc/cpu/cpuregs/_0673_ ;
 wire \soc/cpu/cpuregs/_0674_ ;
 wire \soc/cpu/cpuregs/_0675_ ;
 wire \soc/cpu/cpuregs/_0676_ ;
 wire \soc/cpu/cpuregs/_0677_ ;
 wire \soc/cpu/cpuregs/_0678_ ;
 wire \soc/cpu/cpuregs/_0679_ ;
 wire \soc/cpu/cpuregs/_0680_ ;
 wire \soc/cpu/cpuregs/_0681_ ;
 wire \soc/cpu/cpuregs/_0682_ ;
 wire \soc/cpu/cpuregs/_0683_ ;
 wire \soc/cpu/cpuregs/_0684_ ;
 wire \soc/cpu/cpuregs/_0685_ ;
 wire \soc/cpu/cpuregs/_0686_ ;
 wire \soc/cpu/cpuregs/_0687_ ;
 wire \soc/cpu/cpuregs/_0688_ ;
 wire \soc/cpu/cpuregs/_0689_ ;
 wire \soc/cpu/cpuregs/_0690_ ;
 wire \soc/cpu/cpuregs/_0691_ ;
 wire \soc/cpu/cpuregs/_0692_ ;
 wire \soc/cpu/cpuregs/_0693_ ;
 wire \soc/cpu/cpuregs/_0694_ ;
 wire \soc/cpu/cpuregs/_0695_ ;
 wire \soc/cpu/cpuregs/_0696_ ;
 wire \soc/cpu/cpuregs/_0697_ ;
 wire \soc/cpu/cpuregs/_0698_ ;
 wire \soc/cpu/cpuregs/_0699_ ;
 wire \soc/cpu/cpuregs/_0700_ ;
 wire \soc/cpu/cpuregs/_0701_ ;
 wire \soc/cpu/cpuregs/_0702_ ;
 wire \soc/cpu/cpuregs/_0703_ ;
 wire \soc/cpu/cpuregs/_0704_ ;
 wire \soc/cpu/cpuregs/_0705_ ;
 wire \soc/cpu/cpuregs/_0706_ ;
 wire \soc/cpu/cpuregs/_0707_ ;
 wire \soc/cpu/cpuregs/_0708_ ;
 wire \soc/cpu/cpuregs/_0709_ ;
 wire \soc/cpu/cpuregs/_0710_ ;
 wire \soc/cpu/cpuregs/_0711_ ;
 wire \soc/cpu/cpuregs/_0712_ ;
 wire \soc/cpu/cpuregs/_0713_ ;
 wire \soc/cpu/cpuregs/_0714_ ;
 wire \soc/cpu/cpuregs/_0715_ ;
 wire \soc/cpu/cpuregs/_0716_ ;
 wire \soc/cpu/cpuregs/_0717_ ;
 wire \soc/cpu/cpuregs/_0718_ ;
 wire \soc/cpu/cpuregs/_0719_ ;
 wire \soc/cpu/cpuregs/_0720_ ;
 wire \soc/cpu/cpuregs/_0721_ ;
 wire \soc/cpu/cpuregs/_0722_ ;
 wire \soc/cpu/cpuregs/_0723_ ;
 wire \soc/cpu/cpuregs/_0724_ ;
 wire \soc/cpu/cpuregs/_0725_ ;
 wire \soc/cpu/cpuregs/_0726_ ;
 wire \soc/cpu/cpuregs/_0727_ ;
 wire \soc/cpu/cpuregs/_0728_ ;
 wire \soc/cpu/cpuregs/_0729_ ;
 wire \soc/cpu/cpuregs/_0730_ ;
 wire \soc/cpu/cpuregs/_0731_ ;
 wire \soc/cpu/cpuregs/_0732_ ;
 wire \soc/cpu/cpuregs/_0733_ ;
 wire \soc/cpu/cpuregs/_0734_ ;
 wire \soc/cpu/cpuregs/_0735_ ;
 wire \soc/cpu/cpuregs/_0736_ ;
 wire \soc/cpu/cpuregs/_0737_ ;
 wire \soc/cpu/cpuregs/_0738_ ;
 wire \soc/cpu/cpuregs/_0739_ ;
 wire \soc/cpu/cpuregs/_0740_ ;
 wire \soc/cpu/cpuregs/_0741_ ;
 wire \soc/cpu/cpuregs/_0742_ ;
 wire \soc/cpu/cpuregs/_0743_ ;
 wire \soc/cpu/cpuregs/_0744_ ;
 wire \soc/cpu/cpuregs/_0745_ ;
 wire \soc/cpu/cpuregs/_0746_ ;
 wire \soc/cpu/cpuregs/_0747_ ;
 wire \soc/cpu/cpuregs/_0748_ ;
 wire \soc/cpu/cpuregs/_0749_ ;
 wire \soc/cpu/cpuregs/_0750_ ;
 wire \soc/cpu/cpuregs/_0751_ ;
 wire \soc/cpu/cpuregs/_0752_ ;
 wire \soc/cpu/cpuregs/_0753_ ;
 wire \soc/cpu/cpuregs/_0754_ ;
 wire \soc/cpu/cpuregs/_0755_ ;
 wire \soc/cpu/cpuregs/_0756_ ;
 wire \soc/cpu/cpuregs/_0757_ ;
 wire \soc/cpu/cpuregs/_0758_ ;
 wire \soc/cpu/cpuregs/_0759_ ;
 wire \soc/cpu/cpuregs/_0760_ ;
 wire \soc/cpu/cpuregs/_0761_ ;
 wire \soc/cpu/cpuregs/_0762_ ;
 wire \soc/cpu/cpuregs/_0763_ ;
 wire \soc/cpu/cpuregs/_0764_ ;
 wire \soc/cpu/cpuregs/_0765_ ;
 wire \soc/cpu/cpuregs/_0766_ ;
 wire \soc/cpu/cpuregs/_0767_ ;
 wire \soc/cpu/cpuregs/_0768_ ;
 wire \soc/cpu/cpuregs/_0769_ ;
 wire \soc/cpu/cpuregs/_0770_ ;
 wire \soc/cpu/cpuregs/_0771_ ;
 wire \soc/cpu/cpuregs/_0772_ ;
 wire \soc/cpu/cpuregs/_0773_ ;
 wire \soc/cpu/cpuregs/_0774_ ;
 wire \soc/cpu/cpuregs/_0775_ ;
 wire \soc/cpu/cpuregs/_0776_ ;
 wire \soc/cpu/cpuregs/_0777_ ;
 wire \soc/cpu/cpuregs/_0778_ ;
 wire \soc/cpu/cpuregs/_0779_ ;
 wire \soc/cpu/cpuregs/_0780_ ;
 wire \soc/cpu/cpuregs/_0781_ ;
 wire \soc/cpu/cpuregs/_0782_ ;
 wire \soc/cpu/cpuregs/_0783_ ;
 wire \soc/cpu/cpuregs/_0784_ ;
 wire \soc/cpu/cpuregs/_0785_ ;
 wire \soc/cpu/cpuregs/_0786_ ;
 wire \soc/cpu/cpuregs/_0787_ ;
 wire \soc/cpu/cpuregs/_0788_ ;
 wire \soc/cpu/cpuregs/_0789_ ;
 wire \soc/cpu/cpuregs/_0790_ ;
 wire \soc/cpu/cpuregs/_0791_ ;
 wire \soc/cpu/cpuregs/_0792_ ;
 wire \soc/cpu/cpuregs/_0793_ ;
 wire \soc/cpu/cpuregs/_0794_ ;
 wire \soc/cpu/cpuregs/_0795_ ;
 wire \soc/cpu/cpuregs/_0796_ ;
 wire \soc/cpu/cpuregs/_0797_ ;
 wire \soc/cpu/cpuregs/_0798_ ;
 wire \soc/cpu/cpuregs/_0799_ ;
 wire \soc/cpu/cpuregs/_0800_ ;
 wire \soc/cpu/cpuregs/_0801_ ;
 wire \soc/cpu/cpuregs/_0802_ ;
 wire \soc/cpu/cpuregs/_0803_ ;
 wire \soc/cpu/cpuregs/_0804_ ;
 wire \soc/cpu/cpuregs/_0805_ ;
 wire \soc/cpu/cpuregs/_0806_ ;
 wire \soc/cpu/cpuregs/_0807_ ;
 wire \soc/cpu/cpuregs/_0808_ ;
 wire \soc/cpu/cpuregs/_0809_ ;
 wire \soc/cpu/cpuregs/_0810_ ;
 wire \soc/cpu/cpuregs/_0811_ ;
 wire \soc/cpu/cpuregs/_0812_ ;
 wire \soc/cpu/cpuregs/_0813_ ;
 wire \soc/cpu/cpuregs/_0814_ ;
 wire \soc/cpu/cpuregs/_0815_ ;
 wire \soc/cpu/cpuregs/_0816_ ;
 wire \soc/cpu/cpuregs/_0817_ ;
 wire \soc/cpu/cpuregs/_0818_ ;
 wire \soc/cpu/cpuregs/_0819_ ;
 wire \soc/cpu/cpuregs/_0820_ ;
 wire \soc/cpu/cpuregs/_0821_ ;
 wire \soc/cpu/cpuregs/_0822_ ;
 wire \soc/cpu/cpuregs/_0823_ ;
 wire \soc/cpu/cpuregs/_0824_ ;
 wire \soc/cpu/cpuregs/_0825_ ;
 wire \soc/cpu/cpuregs/_0826_ ;
 wire \soc/cpu/cpuregs/_0827_ ;
 wire \soc/cpu/cpuregs/_0828_ ;
 wire \soc/cpu/cpuregs/_0829_ ;
 wire \soc/cpu/cpuregs/_0830_ ;
 wire \soc/cpu/cpuregs/_0831_ ;
 wire \soc/cpu/cpuregs/_0832_ ;
 wire \soc/cpu/cpuregs/_0833_ ;
 wire \soc/cpu/cpuregs/_0834_ ;
 wire \soc/cpu/cpuregs/_0835_ ;
 wire \soc/cpu/cpuregs/_0836_ ;
 wire \soc/cpu/cpuregs/_0837_ ;
 wire \soc/cpu/cpuregs/_0838_ ;
 wire \soc/cpu/cpuregs/_0839_ ;
 wire \soc/cpu/cpuregs/_0840_ ;
 wire \soc/cpu/cpuregs/_0841_ ;
 wire \soc/cpu/cpuregs/_0842_ ;
 wire \soc/cpu/cpuregs/_0843_ ;
 wire \soc/cpu/cpuregs/_0844_ ;
 wire \soc/cpu/cpuregs/_0845_ ;
 wire \soc/cpu/cpuregs/_0846_ ;
 wire \soc/cpu/cpuregs/_0847_ ;
 wire \soc/cpu/cpuregs/_0848_ ;
 wire \soc/cpu/cpuregs/_0849_ ;
 wire \soc/cpu/cpuregs/_0850_ ;
 wire \soc/cpu/cpuregs/_0851_ ;
 wire \soc/cpu/cpuregs/_0852_ ;
 wire \soc/cpu/cpuregs/_0853_ ;
 wire \soc/cpu/cpuregs/_0854_ ;
 wire \soc/cpu/cpuregs/_0855_ ;
 wire \soc/cpu/cpuregs/_0856_ ;
 wire \soc/cpu/cpuregs/_0857_ ;
 wire \soc/cpu/cpuregs/_0858_ ;
 wire \soc/cpu/cpuregs/_0859_ ;
 wire \soc/cpu/cpuregs/_0860_ ;
 wire \soc/cpu/cpuregs/_0861_ ;
 wire \soc/cpu/cpuregs/_0862_ ;
 wire \soc/cpu/cpuregs/_0863_ ;
 wire \soc/cpu/cpuregs/_0864_ ;
 wire \soc/cpu/cpuregs/_0865_ ;
 wire \soc/cpu/cpuregs/_0866_ ;
 wire \soc/cpu/cpuregs/_0867_ ;
 wire \soc/cpu/cpuregs/_0868_ ;
 wire \soc/cpu/cpuregs/_0869_ ;
 wire \soc/cpu/cpuregs/_0870_ ;
 wire \soc/cpu/cpuregs/_0871_ ;
 wire \soc/cpu/cpuregs/_0872_ ;
 wire \soc/cpu/cpuregs/_0873_ ;
 wire \soc/cpu/cpuregs/_0874_ ;
 wire \soc/cpu/cpuregs/_0875_ ;
 wire \soc/cpu/cpuregs/_0876_ ;
 wire \soc/cpu/cpuregs/_0877_ ;
 wire \soc/cpu/cpuregs/_0878_ ;
 wire \soc/cpu/cpuregs/_0879_ ;
 wire \soc/cpu/cpuregs/_0880_ ;
 wire \soc/cpu/cpuregs/_0881_ ;
 wire \soc/cpu/cpuregs/_0882_ ;
 wire \soc/cpu/cpuregs/_0883_ ;
 wire \soc/cpu/cpuregs/_0884_ ;
 wire \soc/cpu/cpuregs/_0885_ ;
 wire \soc/cpu/cpuregs/_0886_ ;
 wire \soc/cpu/cpuregs/_0887_ ;
 wire \soc/cpu/cpuregs/_0888_ ;
 wire \soc/cpu/cpuregs/_0889_ ;
 wire \soc/cpu/cpuregs/_0890_ ;
 wire \soc/cpu/cpuregs/_0891_ ;
 wire \soc/cpu/cpuregs/_0892_ ;
 wire \soc/cpu/cpuregs/_0893_ ;
 wire \soc/cpu/cpuregs/_0894_ ;
 wire \soc/cpu/cpuregs/_0895_ ;
 wire \soc/cpu/cpuregs/_0896_ ;
 wire \soc/cpu/cpuregs/_0897_ ;
 wire \soc/cpu/cpuregs/_0898_ ;
 wire \soc/cpu/cpuregs/_0899_ ;
 wire \soc/cpu/cpuregs/_0900_ ;
 wire \soc/cpu/cpuregs/_0901_ ;
 wire \soc/cpu/cpuregs/_0902_ ;
 wire \soc/cpu/cpuregs/_0903_ ;
 wire \soc/cpu/cpuregs/_0904_ ;
 wire \soc/cpu/cpuregs/_0905_ ;
 wire \soc/cpu/cpuregs/_0906_ ;
 wire \soc/cpu/cpuregs/_0907_ ;
 wire \soc/cpu/cpuregs/_0908_ ;
 wire \soc/cpu/cpuregs/_0909_ ;
 wire \soc/cpu/cpuregs/_0910_ ;
 wire \soc/cpu/cpuregs/_0911_ ;
 wire \soc/cpu/cpuregs/_0912_ ;
 wire \soc/cpu/cpuregs/_0913_ ;
 wire \soc/cpu/cpuregs/_0914_ ;
 wire \soc/cpu/cpuregs/_0915_ ;
 wire \soc/cpu/cpuregs/_0916_ ;
 wire \soc/cpu/cpuregs/_0917_ ;
 wire \soc/cpu/cpuregs/_0918_ ;
 wire \soc/cpu/cpuregs/_0919_ ;
 wire \soc/cpu/cpuregs/_0920_ ;
 wire \soc/cpu/cpuregs/_0921_ ;
 wire \soc/cpu/cpuregs/_0922_ ;
 wire \soc/cpu/cpuregs/_0923_ ;
 wire \soc/cpu/cpuregs/_0924_ ;
 wire \soc/cpu/cpuregs/_0925_ ;
 wire \soc/cpu/cpuregs/_0926_ ;
 wire \soc/cpu/cpuregs/_0927_ ;
 wire \soc/cpu/cpuregs/_0928_ ;
 wire \soc/cpu/cpuregs/_0929_ ;
 wire \soc/cpu/cpuregs/_0930_ ;
 wire \soc/cpu/cpuregs/_0931_ ;
 wire \soc/cpu/cpuregs/_0932_ ;
 wire \soc/cpu/cpuregs/_0933_ ;
 wire \soc/cpu/cpuregs/_0934_ ;
 wire \soc/cpu/cpuregs/_0935_ ;
 wire \soc/cpu/cpuregs/_0936_ ;
 wire \soc/cpu/cpuregs/_0937_ ;
 wire \soc/cpu/cpuregs/_0938_ ;
 wire \soc/cpu/cpuregs/_0939_ ;
 wire \soc/cpu/cpuregs/_0940_ ;
 wire \soc/cpu/cpuregs/_0941_ ;
 wire \soc/cpu/cpuregs/_0942_ ;
 wire \soc/cpu/cpuregs/_0943_ ;
 wire \soc/cpu/cpuregs/_0944_ ;
 wire \soc/cpu/cpuregs/_0945_ ;
 wire \soc/cpu/cpuregs/_0946_ ;
 wire \soc/cpu/cpuregs/_0947_ ;
 wire \soc/cpu/cpuregs/_0948_ ;
 wire \soc/cpu/cpuregs/_0949_ ;
 wire \soc/cpu/cpuregs/_0950_ ;
 wire \soc/cpu/cpuregs/_0951_ ;
 wire \soc/cpu/cpuregs/_0952_ ;
 wire \soc/cpu/cpuregs/_0953_ ;
 wire \soc/cpu/cpuregs/_0954_ ;
 wire \soc/cpu/cpuregs/_0955_ ;
 wire \soc/cpu/cpuregs/_0956_ ;
 wire \soc/cpu/cpuregs/_0957_ ;
 wire \soc/cpu/cpuregs/_0958_ ;
 wire \soc/cpu/cpuregs/_0959_ ;
 wire \soc/cpu/cpuregs/_0960_ ;
 wire \soc/cpu/cpuregs/_0961_ ;
 wire \soc/cpu/cpuregs/_0962_ ;
 wire \soc/cpu/cpuregs/_0963_ ;
 wire \soc/cpu/cpuregs/_0964_ ;
 wire \soc/cpu/cpuregs/_0965_ ;
 wire \soc/cpu/cpuregs/_0966_ ;
 wire \soc/cpu/cpuregs/_0967_ ;
 wire \soc/cpu/cpuregs/_0968_ ;
 wire \soc/cpu/cpuregs/_0969_ ;
 wire \soc/cpu/cpuregs/_0970_ ;
 wire \soc/cpu/cpuregs/_0971_ ;
 wire \soc/cpu/cpuregs/_0972_ ;
 wire \soc/cpu/cpuregs/_0973_ ;
 wire \soc/cpu/cpuregs/_0974_ ;
 wire \soc/cpu/cpuregs/_0975_ ;
 wire \soc/cpu/cpuregs/_0976_ ;
 wire \soc/cpu/cpuregs/_0977_ ;
 wire \soc/cpu/cpuregs/_0978_ ;
 wire \soc/cpu/cpuregs/_0979_ ;
 wire \soc/cpu/cpuregs/_0980_ ;
 wire \soc/cpu/cpuregs/_0981_ ;
 wire \soc/cpu/cpuregs/_0982_ ;
 wire \soc/cpu/cpuregs/_0983_ ;
 wire \soc/cpu/cpuregs/_0984_ ;
 wire \soc/cpu/cpuregs/_0985_ ;
 wire \soc/cpu/cpuregs/_0986_ ;
 wire \soc/cpu/cpuregs/_0987_ ;
 wire \soc/cpu/cpuregs/_0988_ ;
 wire \soc/cpu/cpuregs/_0989_ ;
 wire \soc/cpu/cpuregs/_0990_ ;
 wire \soc/cpu/cpuregs/_0991_ ;
 wire \soc/cpu/cpuregs/_0992_ ;
 wire \soc/cpu/cpuregs/_0993_ ;
 wire \soc/cpu/cpuregs/_0994_ ;
 wire \soc/cpu/cpuregs/_0995_ ;
 wire \soc/cpu/cpuregs/_0996_ ;
 wire \soc/cpu/cpuregs/_0997_ ;
 wire \soc/cpu/cpuregs/_0998_ ;
 wire \soc/cpu/cpuregs/_0999_ ;
 wire \soc/cpu/cpuregs/_1000_ ;
 wire \soc/cpu/cpuregs/_1001_ ;
 wire \soc/cpu/cpuregs/_1002_ ;
 wire \soc/cpu/cpuregs/_1003_ ;
 wire \soc/cpu/cpuregs/_1004_ ;
 wire \soc/cpu/cpuregs/_1005_ ;
 wire \soc/cpu/cpuregs/_1006_ ;
 wire \soc/cpu/cpuregs/_1007_ ;
 wire \soc/cpu/cpuregs/_1008_ ;
 wire \soc/cpu/cpuregs/_1009_ ;
 wire \soc/cpu/cpuregs/_1010_ ;
 wire \soc/cpu/cpuregs/_1011_ ;
 wire \soc/cpu/cpuregs/_1012_ ;
 wire \soc/cpu/cpuregs/_1013_ ;
 wire \soc/cpu/cpuregs/_1014_ ;
 wire \soc/cpu/cpuregs/_1015_ ;
 wire \soc/cpu/cpuregs/_1016_ ;
 wire \soc/cpu/cpuregs/_1017_ ;
 wire \soc/cpu/cpuregs/_1018_ ;
 wire \soc/cpu/cpuregs/_1019_ ;
 wire \soc/cpu/cpuregs/_1020_ ;
 wire \soc/cpu/cpuregs/_1021_ ;
 wire \soc/cpu/cpuregs/_1022_ ;
 wire \soc/cpu/cpuregs/_1023_ ;
 wire net630;
 wire \soc/cpu/cpuregs/_1025_ ;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire net625;
 wire net624;
 wire net623;
 wire net622;
 wire net621;
 wire \soc/cpu/cpuregs/_1035_ ;
 wire \soc/cpu/cpuregs/_1036_ ;
 wire \soc/cpu/cpuregs/_1037_ ;
 wire net620;
 wire net619;
 wire net618;
 wire net617;
 wire net616;
 wire \soc/cpu/cpuregs/_1043_ ;
 wire net615;
 wire net614;
 wire \soc/cpu/cpuregs/_1046_ ;
 wire net613;
 wire net612;
 wire net611;
 wire net610;
 wire net609;
 wire net608;
 wire \soc/cpu/cpuregs/_1053_ ;
 wire \soc/cpu/cpuregs/_1054_ ;
 wire net607;
 wire net606;
 wire net605;
 wire \soc/cpu/cpuregs/_1058_ ;
 wire \soc/cpu/cpuregs/_1059_ ;
 wire net604;
 wire \soc/cpu/cpuregs/_1061_ ;
 wire \soc/cpu/cpuregs/_1062_ ;
 wire net603;
 wire net602;
 wire net601;
 wire net600;
 wire \soc/cpu/cpuregs/_1067_ ;
 wire \soc/cpu/cpuregs/_1068_ ;
 wire net599;
 wire net598;
 wire net597;
 wire \soc/cpu/cpuregs/_1072_ ;
 wire net596;
 wire \soc/cpu/cpuregs/_1074_ ;
 wire net595;
 wire net594;
 wire net593;
 wire \soc/cpu/cpuregs/_1078_ ;
 wire \soc/cpu/cpuregs/_1079_ ;
 wire net592;
 wire net591;
 wire net590;
 wire \soc/cpu/cpuregs/_1083_ ;
 wire net589;
 wire net588;
 wire \soc/cpu/cpuregs/_1086_ ;
 wire \soc/cpu/cpuregs/_1087_ ;
 wire net587;
 wire \soc/cpu/cpuregs/_1089_ ;
 wire \soc/cpu/cpuregs/_1090_ ;
 wire net586;
 wire \soc/cpu/cpuregs/_1092_ ;
 wire \soc/cpu/cpuregs/_1093_ ;
 wire net585;
 wire net584;
 wire \soc/cpu/cpuregs/_1096_ ;
 wire net583;
 wire \soc/cpu/cpuregs/_1098_ ;
 wire \soc/cpu/cpuregs/_1099_ ;
 wire net582;
 wire \soc/cpu/cpuregs/_1101_ ;
 wire net581;
 wire \soc/cpu/cpuregs/_1103_ ;
 wire \soc/cpu/cpuregs/_1104_ ;
 wire net580;
 wire \soc/cpu/cpuregs/_1106_ ;
 wire net579;
 wire \soc/cpu/cpuregs/_1108_ ;
 wire net578;
 wire net577;
 wire \soc/cpu/cpuregs/_1111_ ;
 wire net576;
 wire net575;
 wire \soc/cpu/cpuregs/_1114_ ;
 wire net574;
 wire \soc/cpu/cpuregs/_1116_ ;
 wire \soc/cpu/cpuregs/_1117_ ;
 wire net573;
 wire \soc/cpu/cpuregs/_1119_ ;
 wire \soc/cpu/cpuregs/_1120_ ;
 wire \soc/cpu/cpuregs/_1121_ ;
 wire net572;
 wire \soc/cpu/cpuregs/_1123_ ;
 wire net571;
 wire net570;
 wire \soc/cpu/cpuregs/_1126_ ;
 wire \soc/cpu/cpuregs/_1127_ ;
 wire net569;
 wire \soc/cpu/cpuregs/_1129_ ;
 wire net568;
 wire \soc/cpu/cpuregs/_1131_ ;
 wire \soc/cpu/cpuregs/_1132_ ;
 wire net567;
 wire \soc/cpu/cpuregs/_1134_ ;
 wire \soc/cpu/cpuregs/_1135_ ;
 wire \soc/cpu/cpuregs/_1136_ ;
 wire \soc/cpu/cpuregs/_1137_ ;
 wire net566;
 wire \soc/cpu/cpuregs/_1139_ ;
 wire \soc/cpu/cpuregs/_1140_ ;
 wire net565;
 wire \soc/cpu/cpuregs/_1142_ ;
 wire \soc/cpu/cpuregs/_1143_ ;
 wire \soc/cpu/cpuregs/_1144_ ;
 wire \soc/cpu/cpuregs/_1145_ ;
 wire \soc/cpu/cpuregs/_1146_ ;
 wire \soc/cpu/cpuregs/_1147_ ;
 wire \soc/cpu/cpuregs/_1148_ ;
 wire \soc/cpu/cpuregs/_1149_ ;
 wire \soc/cpu/cpuregs/_1150_ ;
 wire \soc/cpu/cpuregs/_1151_ ;
 wire \soc/cpu/cpuregs/_1152_ ;
 wire \soc/cpu/cpuregs/_1153_ ;
 wire \soc/cpu/cpuregs/_1154_ ;
 wire \soc/cpu/cpuregs/_1155_ ;
 wire \soc/cpu/cpuregs/_1156_ ;
 wire \soc/cpu/cpuregs/_1157_ ;
 wire \soc/cpu/cpuregs/_1158_ ;
 wire \soc/cpu/cpuregs/_1159_ ;
 wire \soc/cpu/cpuregs/_1160_ ;
 wire \soc/cpu/cpuregs/_1161_ ;
 wire \soc/cpu/cpuregs/_1162_ ;
 wire net564;
 wire net563;
 wire \soc/cpu/cpuregs/_1165_ ;
 wire \soc/cpu/cpuregs/_1166_ ;
 wire net562;
 wire \soc/cpu/cpuregs/_1168_ ;
 wire \soc/cpu/cpuregs/_1169_ ;
 wire \soc/cpu/cpuregs/_1170_ ;
 wire \soc/cpu/cpuregs/_1171_ ;
 wire \soc/cpu/cpuregs/_1172_ ;
 wire \soc/cpu/cpuregs/_1173_ ;
 wire \soc/cpu/cpuregs/_1174_ ;
 wire \soc/cpu/cpuregs/_1175_ ;
 wire net561;
 wire \soc/cpu/cpuregs/_1177_ ;
 wire \soc/cpu/cpuregs/_1178_ ;
 wire \soc/cpu/cpuregs/_1179_ ;
 wire \soc/cpu/cpuregs/_1180_ ;
 wire \soc/cpu/cpuregs/_1181_ ;
 wire net560;
 wire \soc/cpu/cpuregs/_1183_ ;
 wire \soc/cpu/cpuregs/_1184_ ;
 wire \soc/cpu/cpuregs/_1185_ ;
 wire \soc/cpu/cpuregs/_1186_ ;
 wire net559;
 wire \soc/cpu/cpuregs/_1188_ ;
 wire \soc/cpu/cpuregs/_1189_ ;
 wire \soc/cpu/cpuregs/_1190_ ;
 wire \soc/cpu/cpuregs/_1191_ ;
 wire \soc/cpu/cpuregs/_1192_ ;
 wire net558;
 wire \soc/cpu/cpuregs/_1194_ ;
 wire \soc/cpu/cpuregs/_1195_ ;
 wire \soc/cpu/cpuregs/_1196_ ;
 wire \soc/cpu/cpuregs/_1197_ ;
 wire \soc/cpu/cpuregs/_1198_ ;
 wire \soc/cpu/cpuregs/_1199_ ;
 wire \soc/cpu/cpuregs/_1200_ ;
 wire \soc/cpu/cpuregs/_1201_ ;
 wire net557;
 wire \soc/cpu/cpuregs/_1203_ ;
 wire \soc/cpu/cpuregs/_1204_ ;
 wire \soc/cpu/cpuregs/_1205_ ;
 wire net556;
 wire \soc/cpu/cpuregs/_1207_ ;
 wire \soc/cpu/cpuregs/_1208_ ;
 wire net555;
 wire \soc/cpu/cpuregs/_1210_ ;
 wire \soc/cpu/cpuregs/_1211_ ;
 wire net554;
 wire \soc/cpu/cpuregs/_1213_ ;
 wire \soc/cpu/cpuregs/_1214_ ;
 wire \soc/cpu/cpuregs/_1215_ ;
 wire \soc/cpu/cpuregs/_1216_ ;
 wire \soc/cpu/cpuregs/_1217_ ;
 wire \soc/cpu/cpuregs/_1218_ ;
 wire \soc/cpu/cpuregs/_1219_ ;
 wire \soc/cpu/cpuregs/_1220_ ;
 wire \soc/cpu/cpuregs/_1221_ ;
 wire \soc/cpu/cpuregs/_1222_ ;
 wire net553;
 wire \soc/cpu/cpuregs/_1224_ ;
 wire \soc/cpu/cpuregs/_1225_ ;
 wire \soc/cpu/cpuregs/_1226_ ;
 wire \soc/cpu/cpuregs/_1227_ ;
 wire \soc/cpu/cpuregs/_1228_ ;
 wire \soc/cpu/cpuregs/_1229_ ;
 wire \soc/cpu/cpuregs/_1230_ ;
 wire \soc/cpu/cpuregs/_1231_ ;
 wire \soc/cpu/cpuregs/_1232_ ;
 wire \soc/cpu/cpuregs/_1233_ ;
 wire \soc/cpu/cpuregs/_1234_ ;
 wire \soc/cpu/cpuregs/_1235_ ;
 wire \soc/cpu/cpuregs/_1236_ ;
 wire \soc/cpu/cpuregs/_1237_ ;
 wire \soc/cpu/cpuregs/_1238_ ;
 wire \soc/cpu/cpuregs/_1239_ ;
 wire \soc/cpu/cpuregs/_1240_ ;
 wire \soc/cpu/cpuregs/_1241_ ;
 wire net552;
 wire \soc/cpu/cpuregs/_1243_ ;
 wire \soc/cpu/cpuregs/_1244_ ;
 wire net551;
 wire \soc/cpu/cpuregs/_1246_ ;
 wire \soc/cpu/cpuregs/_1247_ ;
 wire \soc/cpu/cpuregs/_1248_ ;
 wire \soc/cpu/cpuregs/_1249_ ;
 wire net550;
 wire net549;
 wire \soc/cpu/cpuregs/_1252_ ;
 wire \soc/cpu/cpuregs/_1253_ ;
 wire \soc/cpu/cpuregs/_1254_ ;
 wire \soc/cpu/cpuregs/_1255_ ;
 wire \soc/cpu/cpuregs/_1256_ ;
 wire \soc/cpu/cpuregs/_1257_ ;
 wire net548;
 wire \soc/cpu/cpuregs/_1259_ ;
 wire \soc/cpu/cpuregs/_1260_ ;
 wire \soc/cpu/cpuregs/_1261_ ;
 wire \soc/cpu/cpuregs/_1262_ ;
 wire \soc/cpu/cpuregs/_1263_ ;
 wire net547;
 wire net546;
 wire \soc/cpu/cpuregs/_1266_ ;
 wire net545;
 wire \soc/cpu/cpuregs/_1268_ ;
 wire \soc/cpu/cpuregs/_1269_ ;
 wire \soc/cpu/cpuregs/_1270_ ;
 wire \soc/cpu/cpuregs/_1271_ ;
 wire \soc/cpu/cpuregs/_1272_ ;
 wire \soc/cpu/cpuregs/_1273_ ;
 wire \soc/cpu/cpuregs/_1274_ ;
 wire \soc/cpu/cpuregs/_1275_ ;
 wire net544;
 wire \soc/cpu/cpuregs/_1277_ ;
 wire \soc/cpu/cpuregs/_1278_ ;
 wire \soc/cpu/cpuregs/_1279_ ;
 wire \soc/cpu/cpuregs/_1280_ ;
 wire \soc/cpu/cpuregs/_1281_ ;
 wire \soc/cpu/cpuregs/_1282_ ;
 wire \soc/cpu/cpuregs/_1283_ ;
 wire \soc/cpu/cpuregs/_1284_ ;
 wire \soc/cpu/cpuregs/_1285_ ;
 wire \soc/cpu/cpuregs/_1286_ ;
 wire \soc/cpu/cpuregs/_1287_ ;
 wire \soc/cpu/cpuregs/_1288_ ;
 wire \soc/cpu/cpuregs/_1289_ ;
 wire \soc/cpu/cpuregs/_1290_ ;
 wire \soc/cpu/cpuregs/_1291_ ;
 wire \soc/cpu/cpuregs/_1292_ ;
 wire \soc/cpu/cpuregs/_1293_ ;
 wire \soc/cpu/cpuregs/_1294_ ;
 wire \soc/cpu/cpuregs/_1295_ ;
 wire \soc/cpu/cpuregs/_1296_ ;
 wire \soc/cpu/cpuregs/_1297_ ;
 wire \soc/cpu/cpuregs/_1298_ ;
 wire \soc/cpu/cpuregs/_1299_ ;
 wire \soc/cpu/cpuregs/_1300_ ;
 wire \soc/cpu/cpuregs/_1301_ ;
 wire \soc/cpu/cpuregs/_1302_ ;
 wire net543;
 wire \soc/cpu/cpuregs/_1304_ ;
 wire \soc/cpu/cpuregs/_1305_ ;
 wire \soc/cpu/cpuregs/_1306_ ;
 wire \soc/cpu/cpuregs/_1307_ ;
 wire \soc/cpu/cpuregs/_1308_ ;
 wire \soc/cpu/cpuregs/_1309_ ;
 wire \soc/cpu/cpuregs/_1310_ ;
 wire net542;
 wire \soc/cpu/cpuregs/_1312_ ;
 wire \soc/cpu/cpuregs/_1313_ ;
 wire \soc/cpu/cpuregs/_1314_ ;
 wire \soc/cpu/cpuregs/_1315_ ;
 wire \soc/cpu/cpuregs/_1316_ ;
 wire \soc/cpu/cpuregs/_1317_ ;
 wire \soc/cpu/cpuregs/_1318_ ;
 wire \soc/cpu/cpuregs/_1319_ ;
 wire \soc/cpu/cpuregs/_1320_ ;
 wire \soc/cpu/cpuregs/_1321_ ;
 wire net541;
 wire \soc/cpu/cpuregs/_1323_ ;
 wire \soc/cpu/cpuregs/_1324_ ;
 wire \soc/cpu/cpuregs/_1325_ ;
 wire \soc/cpu/cpuregs/_1326_ ;
 wire \soc/cpu/cpuregs/_1327_ ;
 wire \soc/cpu/cpuregs/_1328_ ;
 wire \soc/cpu/cpuregs/_1329_ ;
 wire \soc/cpu/cpuregs/_1330_ ;
 wire \soc/cpu/cpuregs/_1331_ ;
 wire \soc/cpu/cpuregs/_1332_ ;
 wire \soc/cpu/cpuregs/_1333_ ;
 wire \soc/cpu/cpuregs/_1334_ ;
 wire \soc/cpu/cpuregs/_1335_ ;
 wire net540;
 wire \soc/cpu/cpuregs/_1337_ ;
 wire \soc/cpu/cpuregs/_1338_ ;
 wire net539;
 wire \soc/cpu/cpuregs/_1340_ ;
 wire \soc/cpu/cpuregs/_1341_ ;
 wire \soc/cpu/cpuregs/_1342_ ;
 wire \soc/cpu/cpuregs/_1343_ ;
 wire \soc/cpu/cpuregs/_1344_ ;
 wire \soc/cpu/cpuregs/_1345_ ;
 wire \soc/cpu/cpuregs/_1346_ ;
 wire \soc/cpu/cpuregs/_1347_ ;
 wire \soc/cpu/cpuregs/_1348_ ;
 wire \soc/cpu/cpuregs/_1349_ ;
 wire net538;
 wire net537;
 wire \soc/cpu/cpuregs/_1352_ ;
 wire \soc/cpu/cpuregs/_1353_ ;
 wire \soc/cpu/cpuregs/_1354_ ;
 wire \soc/cpu/cpuregs/_1355_ ;
 wire \soc/cpu/cpuregs/_1356_ ;
 wire \soc/cpu/cpuregs/_1357_ ;
 wire \soc/cpu/cpuregs/_1358_ ;
 wire \soc/cpu/cpuregs/_1359_ ;
 wire \soc/cpu/cpuregs/_1360_ ;
 wire \soc/cpu/cpuregs/_1361_ ;
 wire \soc/cpu/cpuregs/_1362_ ;
 wire \soc/cpu/cpuregs/_1363_ ;
 wire \soc/cpu/cpuregs/_1364_ ;
 wire \soc/cpu/cpuregs/_1365_ ;
 wire \soc/cpu/cpuregs/_1366_ ;
 wire \soc/cpu/cpuregs/_1367_ ;
 wire \soc/cpu/cpuregs/_1368_ ;
 wire \soc/cpu/cpuregs/_1369_ ;
 wire \soc/cpu/cpuregs/_1370_ ;
 wire \soc/cpu/cpuregs/_1371_ ;
 wire \soc/cpu/cpuregs/_1372_ ;
 wire \soc/cpu/cpuregs/_1373_ ;
 wire \soc/cpu/cpuregs/_1374_ ;
 wire \soc/cpu/cpuregs/_1375_ ;
 wire \soc/cpu/cpuregs/_1376_ ;
 wire \soc/cpu/cpuregs/_1377_ ;
 wire \soc/cpu/cpuregs/_1378_ ;
 wire \soc/cpu/cpuregs/_1379_ ;
 wire \soc/cpu/cpuregs/_1380_ ;
 wire \soc/cpu/cpuregs/_1381_ ;
 wire \soc/cpu/cpuregs/_1382_ ;
 wire \soc/cpu/cpuregs/_1383_ ;
 wire \soc/cpu/cpuregs/_1384_ ;
 wire \soc/cpu/cpuregs/_1385_ ;
 wire \soc/cpu/cpuregs/_1386_ ;
 wire \soc/cpu/cpuregs/_1387_ ;
 wire \soc/cpu/cpuregs/_1388_ ;
 wire \soc/cpu/cpuregs/_1389_ ;
 wire \soc/cpu/cpuregs/_1390_ ;
 wire \soc/cpu/cpuregs/_1391_ ;
 wire \soc/cpu/cpuregs/_1392_ ;
 wire \soc/cpu/cpuregs/_1393_ ;
 wire \soc/cpu/cpuregs/_1394_ ;
 wire \soc/cpu/cpuregs/_1395_ ;
 wire \soc/cpu/cpuregs/_1396_ ;
 wire \soc/cpu/cpuregs/_1397_ ;
 wire \soc/cpu/cpuregs/_1398_ ;
 wire \soc/cpu/cpuregs/_1399_ ;
 wire net536;
 wire \soc/cpu/cpuregs/_1401_ ;
 wire \soc/cpu/cpuregs/_1402_ ;
 wire \soc/cpu/cpuregs/_1403_ ;
 wire \soc/cpu/cpuregs/_1404_ ;
 wire \soc/cpu/cpuregs/_1405_ ;
 wire \soc/cpu/cpuregs/_1406_ ;
 wire \soc/cpu/cpuregs/_1407_ ;
 wire \soc/cpu/cpuregs/_1408_ ;
 wire \soc/cpu/cpuregs/_1409_ ;
 wire net535;
 wire \soc/cpu/cpuregs/_1411_ ;
 wire \soc/cpu/cpuregs/_1412_ ;
 wire \soc/cpu/cpuregs/_1413_ ;
 wire \soc/cpu/cpuregs/_1414_ ;
 wire \soc/cpu/cpuregs/_1415_ ;
 wire \soc/cpu/cpuregs/_1416_ ;
 wire \soc/cpu/cpuregs/_1417_ ;
 wire \soc/cpu/cpuregs/_1418_ ;
 wire net534;
 wire \soc/cpu/cpuregs/_1420_ ;
 wire \soc/cpu/cpuregs/_1421_ ;
 wire \soc/cpu/cpuregs/_1422_ ;
 wire \soc/cpu/cpuregs/_1423_ ;
 wire \soc/cpu/cpuregs/_1424_ ;
 wire \soc/cpu/cpuregs/_1425_ ;
 wire \soc/cpu/cpuregs/_1426_ ;
 wire \soc/cpu/cpuregs/_1427_ ;
 wire \soc/cpu/cpuregs/_1428_ ;
 wire \soc/cpu/cpuregs/_1429_ ;
 wire \soc/cpu/cpuregs/_1430_ ;
 wire \soc/cpu/cpuregs/_1431_ ;
 wire \soc/cpu/cpuregs/_1432_ ;
 wire \soc/cpu/cpuregs/_1433_ ;
 wire \soc/cpu/cpuregs/_1434_ ;
 wire \soc/cpu/cpuregs/_1435_ ;
 wire \soc/cpu/cpuregs/_1436_ ;
 wire \soc/cpu/cpuregs/_1437_ ;
 wire net533;
 wire \soc/cpu/cpuregs/_1439_ ;
 wire \soc/cpu/cpuregs/_1440_ ;
 wire \soc/cpu/cpuregs/_1441_ ;
 wire \soc/cpu/cpuregs/_1442_ ;
 wire net532;
 wire \soc/cpu/cpuregs/_1444_ ;
 wire \soc/cpu/cpuregs/_1445_ ;
 wire \soc/cpu/cpuregs/_1446_ ;
 wire \soc/cpu/cpuregs/_1447_ ;
 wire \soc/cpu/cpuregs/_1448_ ;
 wire net531;
 wire \soc/cpu/cpuregs/_1450_ ;
 wire \soc/cpu/cpuregs/_1451_ ;
 wire \soc/cpu/cpuregs/_1452_ ;
 wire \soc/cpu/cpuregs/_1453_ ;
 wire \soc/cpu/cpuregs/_1454_ ;
 wire \soc/cpu/cpuregs/_1455_ ;
 wire \soc/cpu/cpuregs/_1456_ ;
 wire \soc/cpu/cpuregs/_1457_ ;
 wire \soc/cpu/cpuregs/_1458_ ;
 wire \soc/cpu/cpuregs/_1459_ ;
 wire \soc/cpu/cpuregs/_1460_ ;
 wire \soc/cpu/cpuregs/_1461_ ;
 wire \soc/cpu/cpuregs/_1462_ ;
 wire \soc/cpu/cpuregs/_1463_ ;
 wire \soc/cpu/cpuregs/_1464_ ;
 wire \soc/cpu/cpuregs/_1465_ ;
 wire \soc/cpu/cpuregs/_1466_ ;
 wire \soc/cpu/cpuregs/_1467_ ;
 wire \soc/cpu/cpuregs/_1468_ ;
 wire \soc/cpu/cpuregs/_1469_ ;
 wire \soc/cpu/cpuregs/_1470_ ;
 wire \soc/cpu/cpuregs/_1471_ ;
 wire \soc/cpu/cpuregs/_1472_ ;
 wire \soc/cpu/cpuregs/_1473_ ;
 wire \soc/cpu/cpuregs/_1474_ ;
 wire \soc/cpu/cpuregs/_1475_ ;
 wire \soc/cpu/cpuregs/_1476_ ;
 wire \soc/cpu/cpuregs/_1477_ ;
 wire \soc/cpu/cpuregs/_1478_ ;
 wire \soc/cpu/cpuregs/_1479_ ;
 wire \soc/cpu/cpuregs/_1480_ ;
 wire \soc/cpu/cpuregs/_1481_ ;
 wire \soc/cpu/cpuregs/_1482_ ;
 wire \soc/cpu/cpuregs/_1483_ ;
 wire \soc/cpu/cpuregs/_1484_ ;
 wire \soc/cpu/cpuregs/_1485_ ;
 wire \soc/cpu/cpuregs/_1486_ ;
 wire \soc/cpu/cpuregs/_1487_ ;
 wire \soc/cpu/cpuregs/_1488_ ;
 wire \soc/cpu/cpuregs/_1489_ ;
 wire \soc/cpu/cpuregs/_1490_ ;
 wire \soc/cpu/cpuregs/_1491_ ;
 wire \soc/cpu/cpuregs/_1492_ ;
 wire \soc/cpu/cpuregs/_1493_ ;
 wire \soc/cpu/cpuregs/_1494_ ;
 wire \soc/cpu/cpuregs/_1495_ ;
 wire \soc/cpu/cpuregs/_1496_ ;
 wire \soc/cpu/cpuregs/_1497_ ;
 wire \soc/cpu/cpuregs/_1498_ ;
 wire \soc/cpu/cpuregs/_1499_ ;
 wire \soc/cpu/cpuregs/_1500_ ;
 wire \soc/cpu/cpuregs/_1501_ ;
 wire \soc/cpu/cpuregs/_1502_ ;
 wire \soc/cpu/cpuregs/_1503_ ;
 wire \soc/cpu/cpuregs/_1504_ ;
 wire \soc/cpu/cpuregs/_1505_ ;
 wire \soc/cpu/cpuregs/_1506_ ;
 wire \soc/cpu/cpuregs/_1507_ ;
 wire \soc/cpu/cpuregs/_1508_ ;
 wire \soc/cpu/cpuregs/_1509_ ;
 wire \soc/cpu/cpuregs/_1510_ ;
 wire \soc/cpu/cpuregs/_1511_ ;
 wire \soc/cpu/cpuregs/_1512_ ;
 wire \soc/cpu/cpuregs/_1513_ ;
 wire \soc/cpu/cpuregs/_1514_ ;
 wire \soc/cpu/cpuregs/_1515_ ;
 wire \soc/cpu/cpuregs/_1516_ ;
 wire \soc/cpu/cpuregs/_1517_ ;
 wire \soc/cpu/cpuregs/_1518_ ;
 wire \soc/cpu/cpuregs/_1519_ ;
 wire \soc/cpu/cpuregs/_1520_ ;
 wire \soc/cpu/cpuregs/_1521_ ;
 wire \soc/cpu/cpuregs/_1522_ ;
 wire \soc/cpu/cpuregs/_1523_ ;
 wire \soc/cpu/cpuregs/_1524_ ;
 wire \soc/cpu/cpuregs/_1525_ ;
 wire \soc/cpu/cpuregs/_1526_ ;
 wire \soc/cpu/cpuregs/_1527_ ;
 wire \soc/cpu/cpuregs/_1528_ ;
 wire \soc/cpu/cpuregs/_1529_ ;
 wire \soc/cpu/cpuregs/_1530_ ;
 wire \soc/cpu/cpuregs/_1531_ ;
 wire \soc/cpu/cpuregs/_1532_ ;
 wire \soc/cpu/cpuregs/_1533_ ;
 wire \soc/cpu/cpuregs/_1534_ ;
 wire \soc/cpu/cpuregs/_1535_ ;
 wire \soc/cpu/cpuregs/_1536_ ;
 wire \soc/cpu/cpuregs/_1537_ ;
 wire \soc/cpu/cpuregs/_1538_ ;
 wire \soc/cpu/cpuregs/_1539_ ;
 wire \soc/cpu/cpuregs/_1540_ ;
 wire \soc/cpu/cpuregs/_1541_ ;
 wire \soc/cpu/cpuregs/_1542_ ;
 wire \soc/cpu/cpuregs/_1543_ ;
 wire \soc/cpu/cpuregs/_1544_ ;
 wire \soc/cpu/cpuregs/_1545_ ;
 wire \soc/cpu/cpuregs/_1546_ ;
 wire \soc/cpu/cpuregs/_1547_ ;
 wire \soc/cpu/cpuregs/_1548_ ;
 wire \soc/cpu/cpuregs/_1549_ ;
 wire \soc/cpu/cpuregs/_1550_ ;
 wire \soc/cpu/cpuregs/_1551_ ;
 wire \soc/cpu/cpuregs/_1552_ ;
 wire \soc/cpu/cpuregs/_1553_ ;
 wire \soc/cpu/cpuregs/_1554_ ;
 wire \soc/cpu/cpuregs/_1555_ ;
 wire \soc/cpu/cpuregs/_1556_ ;
 wire \soc/cpu/cpuregs/_1557_ ;
 wire \soc/cpu/cpuregs/_1558_ ;
 wire \soc/cpu/cpuregs/_1559_ ;
 wire \soc/cpu/cpuregs/_1560_ ;
 wire \soc/cpu/cpuregs/_1561_ ;
 wire \soc/cpu/cpuregs/_1562_ ;
 wire \soc/cpu/cpuregs/_1563_ ;
 wire \soc/cpu/cpuregs/_1564_ ;
 wire \soc/cpu/cpuregs/_1565_ ;
 wire \soc/cpu/cpuregs/_1566_ ;
 wire \soc/cpu/cpuregs/_1567_ ;
 wire \soc/cpu/cpuregs/_1568_ ;
 wire \soc/cpu/cpuregs/_1569_ ;
 wire \soc/cpu/cpuregs/_1570_ ;
 wire \soc/cpu/cpuregs/_1571_ ;
 wire \soc/cpu/cpuregs/_1572_ ;
 wire \soc/cpu/cpuregs/_1573_ ;
 wire \soc/cpu/cpuregs/_1574_ ;
 wire \soc/cpu/cpuregs/_1575_ ;
 wire \soc/cpu/cpuregs/_1576_ ;
 wire \soc/cpu/cpuregs/_1577_ ;
 wire \soc/cpu/cpuregs/_1578_ ;
 wire \soc/cpu/cpuregs/_1579_ ;
 wire \soc/cpu/cpuregs/_1580_ ;
 wire \soc/cpu/cpuregs/_1581_ ;
 wire \soc/cpu/cpuregs/_1582_ ;
 wire \soc/cpu/cpuregs/_1583_ ;
 wire \soc/cpu/cpuregs/_1584_ ;
 wire \soc/cpu/cpuregs/_1585_ ;
 wire \soc/cpu/cpuregs/_1586_ ;
 wire \soc/cpu/cpuregs/_1587_ ;
 wire \soc/cpu/cpuregs/_1588_ ;
 wire \soc/cpu/cpuregs/_1589_ ;
 wire \soc/cpu/cpuregs/_1590_ ;
 wire \soc/cpu/cpuregs/_1591_ ;
 wire \soc/cpu/cpuregs/_1592_ ;
 wire \soc/cpu/cpuregs/_1593_ ;
 wire \soc/cpu/cpuregs/_1594_ ;
 wire \soc/cpu/cpuregs/_1595_ ;
 wire \soc/cpu/cpuregs/_1596_ ;
 wire \soc/cpu/cpuregs/_1597_ ;
 wire \soc/cpu/cpuregs/_1598_ ;
 wire \soc/cpu/cpuregs/_1599_ ;
 wire \soc/cpu/cpuregs/_1600_ ;
 wire \soc/cpu/cpuregs/_1601_ ;
 wire \soc/cpu/cpuregs/_1602_ ;
 wire \soc/cpu/cpuregs/_1603_ ;
 wire \soc/cpu/cpuregs/_1604_ ;
 wire \soc/cpu/cpuregs/_1605_ ;
 wire \soc/cpu/cpuregs/_1606_ ;
 wire \soc/cpu/cpuregs/_1607_ ;
 wire \soc/cpu/cpuregs/_1608_ ;
 wire \soc/cpu/cpuregs/_1609_ ;
 wire \soc/cpu/cpuregs/_1610_ ;
 wire \soc/cpu/cpuregs/_1611_ ;
 wire \soc/cpu/cpuregs/_1612_ ;
 wire \soc/cpu/cpuregs/_1613_ ;
 wire \soc/cpu/cpuregs/_1614_ ;
 wire \soc/cpu/cpuregs/_1615_ ;
 wire \soc/cpu/cpuregs/_1616_ ;
 wire \soc/cpu/cpuregs/_1617_ ;
 wire \soc/cpu/cpuregs/_1618_ ;
 wire \soc/cpu/cpuregs/_1619_ ;
 wire \soc/cpu/cpuregs/_1620_ ;
 wire \soc/cpu/cpuregs/_1621_ ;
 wire \soc/cpu/cpuregs/_1622_ ;
 wire \soc/cpu/cpuregs/_1623_ ;
 wire \soc/cpu/cpuregs/_1624_ ;
 wire \soc/cpu/cpuregs/_1625_ ;
 wire \soc/cpu/cpuregs/_1626_ ;
 wire \soc/cpu/cpuregs/_1627_ ;
 wire \soc/cpu/cpuregs/_1628_ ;
 wire \soc/cpu/cpuregs/_1629_ ;
 wire \soc/cpu/cpuregs/_1630_ ;
 wire \soc/cpu/cpuregs/_1631_ ;
 wire \soc/cpu/cpuregs/_1632_ ;
 wire \soc/cpu/cpuregs/_1633_ ;
 wire \soc/cpu/cpuregs/_1634_ ;
 wire \soc/cpu/cpuregs/_1635_ ;
 wire \soc/cpu/cpuregs/_1636_ ;
 wire \soc/cpu/cpuregs/_1637_ ;
 wire \soc/cpu/cpuregs/_1638_ ;
 wire \soc/cpu/cpuregs/_1639_ ;
 wire \soc/cpu/cpuregs/_1640_ ;
 wire \soc/cpu/cpuregs/_1641_ ;
 wire \soc/cpu/cpuregs/_1642_ ;
 wire \soc/cpu/cpuregs/_1643_ ;
 wire \soc/cpu/cpuregs/_1644_ ;
 wire \soc/cpu/cpuregs/_1645_ ;
 wire \soc/cpu/cpuregs/_1646_ ;
 wire \soc/cpu/cpuregs/_1647_ ;
 wire \soc/cpu/cpuregs/_1648_ ;
 wire \soc/cpu/cpuregs/_1649_ ;
 wire \soc/cpu/cpuregs/_1650_ ;
 wire \soc/cpu/cpuregs/_1651_ ;
 wire \soc/cpu/cpuregs/_1652_ ;
 wire \soc/cpu/cpuregs/_1653_ ;
 wire \soc/cpu/cpuregs/_1654_ ;
 wire \soc/cpu/cpuregs/_1655_ ;
 wire \soc/cpu/cpuregs/_1656_ ;
 wire \soc/cpu/cpuregs/_1657_ ;
 wire \soc/cpu/cpuregs/_1658_ ;
 wire \soc/cpu/cpuregs/_1659_ ;
 wire \soc/cpu/cpuregs/_1660_ ;
 wire \soc/cpu/cpuregs/_1661_ ;
 wire \soc/cpu/cpuregs/_1662_ ;
 wire \soc/cpu/cpuregs/_1663_ ;
 wire net530;
 wire net529;
 wire net528;
 wire net527;
 wire net526;
 wire net525;
 wire net524;
 wire net523;
 wire net522;
 wire net521;
 wire net520;
 wire \soc/cpu/cpuregs/_1675_ ;
 wire \soc/cpu/cpuregs/_1676_ ;
 wire \soc/cpu/cpuregs/_1677_ ;
 wire net519;
 wire net518;
 wire net517;
 wire net516;
 wire net515;
 wire \soc/cpu/cpuregs/_1683_ ;
 wire net514;
 wire net513;
 wire \soc/cpu/cpuregs/_1686_ ;
 wire net512;
 wire net511;
 wire net510;
 wire net509;
 wire net508;
 wire \soc/cpu/cpuregs/_1692_ ;
 wire \soc/cpu/cpuregs/_1693_ ;
 wire net507;
 wire net506;
 wire net505;
 wire net504;
 wire \soc/cpu/cpuregs/_1698_ ;
 wire \soc/cpu/cpuregs/_1699_ ;
 wire net503;
 wire net502;
 wire \soc/cpu/cpuregs/_1702_ ;
 wire \soc/cpu/cpuregs/_1703_ ;
 wire net501;
 wire net500;
 wire net499;
 wire net498;
 wire \soc/cpu/cpuregs/_1708_ ;
 wire \soc/cpu/cpuregs/_1709_ ;
 wire net497;
 wire net496;
 wire net495;
 wire \soc/cpu/cpuregs/_1713_ ;
 wire net494;
 wire \soc/cpu/cpuregs/_1715_ ;
 wire net493;
 wire net492;
 wire clknet_3_7_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_5_0_clk;
 wire \soc/cpu/cpuregs/_1721_ ;
 wire \soc/cpu/cpuregs/_1722_ ;
 wire clknet_3_4_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_1_0_clk;
 wire \soc/cpu/cpuregs/_1727_ ;
 wire clknet_3_0_0_clk;
 wire \soc/cpu/cpuregs/_1729_ ;
 wire clknet_2_3_0_clk;
 wire clknet_2_2_0_clk;
 wire \soc/cpu/cpuregs/_1732_ ;
 wire clknet_2_1_0_clk;
 wire \soc/cpu/cpuregs/_1734_ ;
 wire clknet_2_0_0_clk;
 wire \soc/cpu/cpuregs/_1736_ ;
 wire clknet_1_1_1_clk;
 wire \soc/cpu/cpuregs/_1738_ ;
 wire clknet_1_1_0_clk;
 wire clknet_1_0_1_clk;
 wire \soc/cpu/cpuregs/_1741_ ;
 wire \soc/cpu/cpuregs/_1742_ ;
 wire \soc/cpu/cpuregs/_1743_ ;
 wire clknet_1_0_0_clk;
 wire \soc/cpu/cpuregs/_1745_ ;
 wire \soc/cpu/cpuregs/_1746_ ;
 wire \soc/cpu/cpuregs/_1747_ ;
 wire \soc/cpu/cpuregs/_1748_ ;
 wire \soc/cpu/cpuregs/_1749_ ;
 wire \soc/cpu/cpuregs/_1750_ ;
 wire \soc/cpu/cpuregs/_1751_ ;
 wire \soc/cpu/cpuregs/_1752_ ;
 wire \soc/cpu/cpuregs/_1753_ ;
 wire \soc/cpu/cpuregs/_1754_ ;
 wire clknet_0_clk;
 wire \soc/cpu/cpuregs/_1756_ ;
 wire \soc/cpu/cpuregs/_1757_ ;
 wire \soc/cpu/cpuregs/_1758_ ;
 wire \soc/cpu/cpuregs/_1759_ ;
 wire \soc/cpu/cpuregs/_1760_ ;
 wire clknet_leaf_94_clk;
 wire \soc/cpu/cpuregs/_1762_ ;
 wire \soc/cpu/cpuregs/_1763_ ;
 wire \soc/cpu/cpuregs/_1764_ ;
 wire \soc/cpu/cpuregs/_1765_ ;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_92_clk;
 wire \soc/cpu/cpuregs/_1768_ ;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_90_clk;
 wire \soc/cpu/cpuregs/_1771_ ;
 wire clknet_leaf_89_clk;
 wire \soc/cpu/cpuregs/_1773_ ;
 wire clknet_leaf_88_clk;
 wire \soc/cpu/cpuregs/_1775_ ;
 wire \soc/cpu/cpuregs/_1776_ ;
 wire \soc/cpu/cpuregs/_1777_ ;
 wire \soc/cpu/cpuregs/_1778_ ;
 wire \soc/cpu/cpuregs/_1779_ ;
 wire \soc/cpu/cpuregs/_1780_ ;
 wire \soc/cpu/cpuregs/_1781_ ;
 wire clknet_leaf_87_clk;
 wire \soc/cpu/cpuregs/_1783_ ;
 wire \soc/cpu/cpuregs/_1784_ ;
 wire \soc/cpu/cpuregs/_1785_ ;
 wire \soc/cpu/cpuregs/_1786_ ;
 wire \soc/cpu/cpuregs/_1787_ ;
 wire \soc/cpu/cpuregs/_1788_ ;
 wire \soc/cpu/cpuregs/_1789_ ;
 wire \soc/cpu/cpuregs/_1790_ ;
 wire clknet_leaf_86_clk;
 wire \soc/cpu/cpuregs/_1792_ ;
 wire \soc/cpu/cpuregs/_1793_ ;
 wire \soc/cpu/cpuregs/_1794_ ;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_84_clk;
 wire \soc/cpu/cpuregs/_1797_ ;
 wire \soc/cpu/cpuregs/_1798_ ;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_82_clk;
 wire \soc/cpu/cpuregs/_1801_ ;
 wire \soc/cpu/cpuregs/_1802_ ;
 wire \soc/cpu/cpuregs/_1803_ ;
 wire \soc/cpu/cpuregs/_1804_ ;
 wire \soc/cpu/cpuregs/_1805_ ;
 wire \soc/cpu/cpuregs/_1806_ ;
 wire \soc/cpu/cpuregs/_1807_ ;
 wire \soc/cpu/cpuregs/_1808_ ;
 wire \soc/cpu/cpuregs/_1809_ ;
 wire \soc/cpu/cpuregs/_1810_ ;
 wire clknet_leaf_81_clk;
 wire \soc/cpu/cpuregs/_1812_ ;
 wire \soc/cpu/cpuregs/_1813_ ;
 wire \soc/cpu/cpuregs/_1814_ ;
 wire \soc/cpu/cpuregs/_1815_ ;
 wire clknet_leaf_80_clk;
 wire \soc/cpu/cpuregs/_1817_ ;
 wire \soc/cpu/cpuregs/_1818_ ;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_77_clk;
 wire \soc/cpu/cpuregs/_1822_ ;
 wire \soc/cpu/cpuregs/_1823_ ;
 wire \soc/cpu/cpuregs/_1824_ ;
 wire \soc/cpu/cpuregs/_1825_ ;
 wire \soc/cpu/cpuregs/_1826_ ;
 wire \soc/cpu/cpuregs/_1827_ ;
 wire \soc/cpu/cpuregs/_1828_ ;
 wire \soc/cpu/cpuregs/_1829_ ;
 wire clknet_leaf_76_clk;
 wire \soc/cpu/cpuregs/_1831_ ;
 wire \soc/cpu/cpuregs/_1832_ ;
 wire \soc/cpu/cpuregs/_1833_ ;
 wire \soc/cpu/cpuregs/_1834_ ;
 wire \soc/cpu/cpuregs/_1835_ ;
 wire \soc/cpu/cpuregs/_1836_ ;
 wire \soc/cpu/cpuregs/_1837_ ;
 wire \soc/cpu/cpuregs/_1838_ ;
 wire \soc/cpu/cpuregs/_1839_ ;
 wire \soc/cpu/cpuregs/_1840_ ;
 wire \soc/cpu/cpuregs/_1841_ ;
 wire clknet_leaf_75_clk;
 wire \soc/cpu/cpuregs/_1843_ ;
 wire \soc/cpu/cpuregs/_1844_ ;
 wire \soc/cpu/cpuregs/_1845_ ;
 wire \soc/cpu/cpuregs/_1846_ ;
 wire \soc/cpu/cpuregs/_1847_ ;
 wire clknet_leaf_74_clk;
 wire \soc/cpu/cpuregs/_1849_ ;
 wire \soc/cpu/cpuregs/_1850_ ;
 wire \soc/cpu/cpuregs/_1851_ ;
 wire \soc/cpu/cpuregs/_1852_ ;
 wire \soc/cpu/cpuregs/_1853_ ;
 wire \soc/cpu/cpuregs/_1854_ ;
 wire \soc/cpu/cpuregs/_1855_ ;
 wire \soc/cpu/cpuregs/_1856_ ;
 wire \soc/cpu/cpuregs/_1857_ ;
 wire \soc/cpu/cpuregs/_1858_ ;
 wire \soc/cpu/cpuregs/_1859_ ;
 wire \soc/cpu/cpuregs/_1860_ ;
 wire \soc/cpu/cpuregs/_1861_ ;
 wire \soc/cpu/cpuregs/_1862_ ;
 wire \soc/cpu/cpuregs/_1863_ ;
 wire \soc/cpu/cpuregs/_1864_ ;
 wire \soc/cpu/cpuregs/_1865_ ;
 wire clknet_leaf_73_clk;
 wire \soc/cpu/cpuregs/_1867_ ;
 wire clknet_leaf_72_clk;
 wire \soc/cpu/cpuregs/_1869_ ;
 wire clknet_leaf_71_clk;
 wire \soc/cpu/cpuregs/_1871_ ;
 wire \soc/cpu/cpuregs/_1872_ ;
 wire \soc/cpu/cpuregs/_1873_ ;
 wire \soc/cpu/cpuregs/_1874_ ;
 wire \soc/cpu/cpuregs/_1875_ ;
 wire \soc/cpu/cpuregs/_1876_ ;
 wire \soc/cpu/cpuregs/_1877_ ;
 wire \soc/cpu/cpuregs/_1878_ ;
 wire \soc/cpu/cpuregs/_1879_ ;
 wire \soc/cpu/cpuregs/_1880_ ;
 wire \soc/cpu/cpuregs/_1881_ ;
 wire \soc/cpu/cpuregs/_1882_ ;
 wire \soc/cpu/cpuregs/_1883_ ;
 wire \soc/cpu/cpuregs/_1884_ ;
 wire \soc/cpu/cpuregs/_1885_ ;
 wire \soc/cpu/cpuregs/_1886_ ;
 wire \soc/cpu/cpuregs/_1887_ ;
 wire \soc/cpu/cpuregs/_1888_ ;
 wire \soc/cpu/cpuregs/_1889_ ;
 wire \soc/cpu/cpuregs/_1890_ ;
 wire clknet_leaf_70_clk;
 wire \soc/cpu/cpuregs/_1892_ ;
 wire \soc/cpu/cpuregs/_1893_ ;
 wire \soc/cpu/cpuregs/_1894_ ;
 wire \soc/cpu/cpuregs/_1895_ ;
 wire \soc/cpu/cpuregs/_1896_ ;
 wire clknet_leaf_69_clk;
 wire \soc/cpu/cpuregs/_1898_ ;
 wire \soc/cpu/cpuregs/_1899_ ;
 wire clknet_leaf_68_clk;
 wire \soc/cpu/cpuregs/_1901_ ;
 wire \soc/cpu/cpuregs/_1902_ ;
 wire \soc/cpu/cpuregs/_1903_ ;
 wire \soc/cpu/cpuregs/_1904_ ;
 wire \soc/cpu/cpuregs/_1905_ ;
 wire \soc/cpu/cpuregs/_1906_ ;
 wire \soc/cpu/cpuregs/_1907_ ;
 wire \soc/cpu/cpuregs/_1908_ ;
 wire \soc/cpu/cpuregs/_1909_ ;
 wire \soc/cpu/cpuregs/_1910_ ;
 wire \soc/cpu/cpuregs/_1911_ ;
 wire clknet_leaf_67_clk;
 wire \soc/cpu/cpuregs/_1913_ ;
 wire \soc/cpu/cpuregs/_1914_ ;
 wire \soc/cpu/cpuregs/_1915_ ;
 wire \soc/cpu/cpuregs/_1916_ ;
 wire \soc/cpu/cpuregs/_1917_ ;
 wire clknet_leaf_66_clk;
 wire \soc/cpu/cpuregs/_1919_ ;
 wire \soc/cpu/cpuregs/_1920_ ;
 wire \soc/cpu/cpuregs/_1921_ ;
 wire \soc/cpu/cpuregs/_1922_ ;
 wire \soc/cpu/cpuregs/_1923_ ;
 wire \soc/cpu/cpuregs/_1924_ ;
 wire \soc/cpu/cpuregs/_1925_ ;
 wire clknet_leaf_65_clk;
 wire \soc/cpu/cpuregs/_1927_ ;
 wire clknet_leaf_63_clk;
 wire \soc/cpu/cpuregs/_1929_ ;
 wire \soc/cpu/cpuregs/_1930_ ;
 wire \soc/cpu/cpuregs/_1931_ ;
 wire \soc/cpu/cpuregs/_1932_ ;
 wire \soc/cpu/cpuregs/_1933_ ;
 wire \soc/cpu/cpuregs/_1934_ ;
 wire clknet_leaf_62_clk;
 wire \soc/cpu/cpuregs/_1936_ ;
 wire \soc/cpu/cpuregs/_1937_ ;
 wire \soc/cpu/cpuregs/_1938_ ;
 wire \soc/cpu/cpuregs/_1939_ ;
 wire \soc/cpu/cpuregs/_1940_ ;
 wire \soc/cpu/cpuregs/_1941_ ;
 wire \soc/cpu/cpuregs/_1942_ ;
 wire \soc/cpu/cpuregs/_1943_ ;
 wire \soc/cpu/cpuregs/_1944_ ;
 wire \soc/cpu/cpuregs/_1945_ ;
 wire \soc/cpu/cpuregs/_1946_ ;
 wire \soc/cpu/cpuregs/_1947_ ;
 wire \soc/cpu/cpuregs/_1948_ ;
 wire \soc/cpu/cpuregs/_1949_ ;
 wire \soc/cpu/cpuregs/_1950_ ;
 wire \soc/cpu/cpuregs/_1951_ ;
 wire \soc/cpu/cpuregs/_1952_ ;
 wire \soc/cpu/cpuregs/_1953_ ;
 wire \soc/cpu/cpuregs/_1954_ ;
 wire \soc/cpu/cpuregs/_1955_ ;
 wire \soc/cpu/cpuregs/_1956_ ;
 wire \soc/cpu/cpuregs/_1957_ ;
 wire \soc/cpu/cpuregs/_1958_ ;
 wire \soc/cpu/cpuregs/_1959_ ;
 wire \soc/cpu/cpuregs/_1960_ ;
 wire \soc/cpu/cpuregs/_1961_ ;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_60_clk;
 wire \soc/cpu/cpuregs/_1964_ ;
 wire \soc/cpu/cpuregs/_1965_ ;
 wire \soc/cpu/cpuregs/_1966_ ;
 wire \soc/cpu/cpuregs/_1967_ ;
 wire \soc/cpu/cpuregs/_1968_ ;
 wire \soc/cpu/cpuregs/_1969_ ;
 wire \soc/cpu/cpuregs/_1970_ ;
 wire \soc/cpu/cpuregs/_1971_ ;
 wire \soc/cpu/cpuregs/_1972_ ;
 wire \soc/cpu/cpuregs/_1973_ ;
 wire \soc/cpu/cpuregs/_1974_ ;
 wire \soc/cpu/cpuregs/_1975_ ;
 wire \soc/cpu/cpuregs/_1976_ ;
 wire clknet_leaf_59_clk;
 wire \soc/cpu/cpuregs/_1978_ ;
 wire \soc/cpu/cpuregs/_1979_ ;
 wire clknet_leaf_58_clk;
 wire \soc/cpu/cpuregs/_1981_ ;
 wire \soc/cpu/cpuregs/_1982_ ;
 wire \soc/cpu/cpuregs/_1983_ ;
 wire clknet_leaf_57_clk;
 wire \soc/cpu/cpuregs/_1985_ ;
 wire \soc/cpu/cpuregs/_1986_ ;
 wire \soc/cpu/cpuregs/_1987_ ;
 wire \soc/cpu/cpuregs/_1988_ ;
 wire \soc/cpu/cpuregs/_1989_ ;
 wire \soc/cpu/cpuregs/_1990_ ;
 wire \soc/cpu/cpuregs/_1991_ ;
 wire \soc/cpu/cpuregs/_1992_ ;
 wire \soc/cpu/cpuregs/_1993_ ;
 wire \soc/cpu/cpuregs/_1994_ ;
 wire \soc/cpu/cpuregs/_1995_ ;
 wire \soc/cpu/cpuregs/_1996_ ;
 wire \soc/cpu/cpuregs/_1997_ ;
 wire \soc/cpu/cpuregs/_1998_ ;
 wire \soc/cpu/cpuregs/_1999_ ;
 wire \soc/cpu/cpuregs/_2000_ ;
 wire \soc/cpu/cpuregs/_2001_ ;
 wire \soc/cpu/cpuregs/_2002_ ;
 wire \soc/cpu/cpuregs/_2003_ ;
 wire \soc/cpu/cpuregs/_2004_ ;
 wire \soc/cpu/cpuregs/_2005_ ;
 wire \soc/cpu/cpuregs/_2006_ ;
 wire \soc/cpu/cpuregs/_2007_ ;
 wire \soc/cpu/cpuregs/_2008_ ;
 wire \soc/cpu/cpuregs/_2009_ ;
 wire \soc/cpu/cpuregs/_2010_ ;
 wire \soc/cpu/cpuregs/_2011_ ;
 wire \soc/cpu/cpuregs/_2012_ ;
 wire \soc/cpu/cpuregs/_2013_ ;
 wire \soc/cpu/cpuregs/_2014_ ;
 wire \soc/cpu/cpuregs/_2015_ ;
 wire \soc/cpu/cpuregs/_2016_ ;
 wire \soc/cpu/cpuregs/_2017_ ;
 wire \soc/cpu/cpuregs/_2018_ ;
 wire \soc/cpu/cpuregs/_2019_ ;
 wire \soc/cpu/cpuregs/_2020_ ;
 wire \soc/cpu/cpuregs/_2021_ ;
 wire \soc/cpu/cpuregs/_2022_ ;
 wire \soc/cpu/cpuregs/_2023_ ;
 wire \soc/cpu/cpuregs/_2024_ ;
 wire \soc/cpu/cpuregs/_2025_ ;
 wire \soc/cpu/cpuregs/_2026_ ;
 wire \soc/cpu/cpuregs/_2027_ ;
 wire \soc/cpu/cpuregs/_2028_ ;
 wire \soc/cpu/cpuregs/_2029_ ;
 wire \soc/cpu/cpuregs/_2030_ ;
 wire \soc/cpu/cpuregs/_2031_ ;
 wire \soc/cpu/cpuregs/_2032_ ;
 wire \soc/cpu/cpuregs/_2033_ ;
 wire \soc/cpu/cpuregs/_2034_ ;
 wire \soc/cpu/cpuregs/_2035_ ;
 wire \soc/cpu/cpuregs/_2036_ ;
 wire \soc/cpu/cpuregs/_2037_ ;
 wire \soc/cpu/cpuregs/_2038_ ;
 wire \soc/cpu/cpuregs/_2039_ ;
 wire \soc/cpu/cpuregs/_2040_ ;
 wire \soc/cpu/cpuregs/_2041_ ;
 wire \soc/cpu/cpuregs/_2042_ ;
 wire clknet_leaf_56_clk;
 wire \soc/cpu/cpuregs/_2044_ ;
 wire \soc/cpu/cpuregs/_2045_ ;
 wire \soc/cpu/cpuregs/_2046_ ;
 wire \soc/cpu/cpuregs/_2047_ ;
 wire \soc/cpu/cpuregs/_2048_ ;
 wire \soc/cpu/cpuregs/_2049_ ;
 wire \soc/cpu/cpuregs/_2050_ ;
 wire \soc/cpu/cpuregs/_2051_ ;
 wire \soc/cpu/cpuregs/_2052_ ;
 wire \soc/cpu/cpuregs/_2053_ ;
 wire \soc/cpu/cpuregs/_2054_ ;
 wire \soc/cpu/cpuregs/_2055_ ;
 wire \soc/cpu/cpuregs/_2056_ ;
 wire \soc/cpu/cpuregs/_2057_ ;
 wire \soc/cpu/cpuregs/_2058_ ;
 wire \soc/cpu/cpuregs/_2059_ ;
 wire \soc/cpu/cpuregs/_2060_ ;
 wire \soc/cpu/cpuregs/_2061_ ;
 wire \soc/cpu/cpuregs/_2062_ ;
 wire \soc/cpu/cpuregs/_2063_ ;
 wire clknet_leaf_55_clk;
 wire \soc/cpu/cpuregs/_2065_ ;
 wire \soc/cpu/cpuregs/_2066_ ;
 wire \soc/cpu/cpuregs/_2067_ ;
 wire \soc/cpu/cpuregs/_2068_ ;
 wire \soc/cpu/cpuregs/_2069_ ;
 wire \soc/cpu/cpuregs/_2070_ ;
 wire \soc/cpu/cpuregs/_2071_ ;
 wire \soc/cpu/cpuregs/_2072_ ;
 wire \soc/cpu/cpuregs/_2073_ ;
 wire \soc/cpu/cpuregs/_2074_ ;
 wire \soc/cpu/cpuregs/_2075_ ;
 wire \soc/cpu/cpuregs/_2076_ ;
 wire \soc/cpu/cpuregs/_2077_ ;
 wire \soc/cpu/cpuregs/_2078_ ;
 wire \soc/cpu/cpuregs/_2079_ ;
 wire \soc/cpu/cpuregs/_2080_ ;
 wire \soc/cpu/cpuregs/_2081_ ;
 wire \soc/cpu/cpuregs/_2082_ ;
 wire \soc/cpu/cpuregs/_2083_ ;
 wire \soc/cpu/cpuregs/_2084_ ;
 wire \soc/cpu/cpuregs/_2085_ ;
 wire \soc/cpu/cpuregs/_2086_ ;
 wire \soc/cpu/cpuregs/_2087_ ;
 wire \soc/cpu/cpuregs/_2088_ ;
 wire \soc/cpu/cpuregs/_2089_ ;
 wire clknet_leaf_54_clk;
 wire \soc/cpu/cpuregs/_2091_ ;
 wire \soc/cpu/cpuregs/_2092_ ;
 wire \soc/cpu/cpuregs/_2093_ ;
 wire \soc/cpu/cpuregs/_2094_ ;
 wire \soc/cpu/cpuregs/_2095_ ;
 wire \soc/cpu/cpuregs/_2096_ ;
 wire \soc/cpu/cpuregs/_2097_ ;
 wire \soc/cpu/cpuregs/_2098_ ;
 wire \soc/cpu/cpuregs/_2099_ ;
 wire \soc/cpu/cpuregs/_2100_ ;
 wire \soc/cpu/cpuregs/_2101_ ;
 wire \soc/cpu/cpuregs/_2102_ ;
 wire \soc/cpu/cpuregs/_2103_ ;
 wire \soc/cpu/cpuregs/_2104_ ;
 wire \soc/cpu/cpuregs/_2105_ ;
 wire \soc/cpu/cpuregs/_2106_ ;
 wire \soc/cpu/cpuregs/_2107_ ;
 wire \soc/cpu/cpuregs/_2108_ ;
 wire \soc/cpu/cpuregs/_2109_ ;
 wire \soc/cpu/cpuregs/_2110_ ;
 wire \soc/cpu/cpuregs/_2111_ ;
 wire \soc/cpu/cpuregs/_2112_ ;
 wire \soc/cpu/cpuregs/_2113_ ;
 wire \soc/cpu/cpuregs/_2114_ ;
 wire \soc/cpu/cpuregs/_2115_ ;
 wire \soc/cpu/cpuregs/_2116_ ;
 wire \soc/cpu/cpuregs/_2117_ ;
 wire \soc/cpu/cpuregs/_2118_ ;
 wire \soc/cpu/cpuregs/_2119_ ;
 wire \soc/cpu/cpuregs/_2120_ ;
 wire \soc/cpu/cpuregs/_2121_ ;
 wire \soc/cpu/cpuregs/_2122_ ;
 wire \soc/cpu/cpuregs/_2123_ ;
 wire \soc/cpu/cpuregs/_2124_ ;
 wire \soc/cpu/cpuregs/_2125_ ;
 wire \soc/cpu/cpuregs/_2126_ ;
 wire \soc/cpu/cpuregs/_2127_ ;
 wire \soc/cpu/cpuregs/_2128_ ;
 wire \soc/cpu/cpuregs/_2129_ ;
 wire \soc/cpu/cpuregs/_2130_ ;
 wire \soc/cpu/cpuregs/_2131_ ;
 wire \soc/cpu/cpuregs/_2132_ ;
 wire \soc/cpu/cpuregs/_2133_ ;
 wire \soc/cpu/cpuregs/_2134_ ;
 wire \soc/cpu/cpuregs/_2135_ ;
 wire \soc/cpu/cpuregs/_2136_ ;
 wire \soc/cpu/cpuregs/_2137_ ;
 wire \soc/cpu/cpuregs/_2138_ ;
 wire \soc/cpu/cpuregs/_2139_ ;
 wire \soc/cpu/cpuregs/_2140_ ;
 wire \soc/cpu/cpuregs/_2141_ ;
 wire \soc/cpu/cpuregs/_2142_ ;
 wire \soc/cpu/cpuregs/_2143_ ;
 wire \soc/cpu/cpuregs/_2144_ ;
 wire \soc/cpu/cpuregs/_2145_ ;
 wire \soc/cpu/cpuregs/_2146_ ;
 wire \soc/cpu/cpuregs/_2147_ ;
 wire \soc/cpu/cpuregs/_2148_ ;
 wire \soc/cpu/cpuregs/_2149_ ;
 wire \soc/cpu/cpuregs/_2150_ ;
 wire \soc/cpu/cpuregs/_2151_ ;
 wire \soc/cpu/cpuregs/_2152_ ;
 wire \soc/cpu/cpuregs/_2153_ ;
 wire \soc/cpu/cpuregs/_2154_ ;
 wire \soc/cpu/cpuregs/_2155_ ;
 wire \soc/cpu/cpuregs/_2156_ ;
 wire \soc/cpu/cpuregs/_2157_ ;
 wire \soc/cpu/cpuregs/_2158_ ;
 wire \soc/cpu/cpuregs/_2159_ ;
 wire \soc/cpu/cpuregs/_2160_ ;
 wire \soc/cpu/cpuregs/_2161_ ;
 wire \soc/cpu/cpuregs/_2162_ ;
 wire \soc/cpu/cpuregs/_2163_ ;
 wire \soc/cpu/cpuregs/_2164_ ;
 wire \soc/cpu/cpuregs/_2165_ ;
 wire \soc/cpu/cpuregs/_2166_ ;
 wire \soc/cpu/cpuregs/_2167_ ;
 wire \soc/cpu/cpuregs/_2168_ ;
 wire \soc/cpu/cpuregs/_2169_ ;
 wire \soc/cpu/cpuregs/_2170_ ;
 wire \soc/cpu/cpuregs/_2171_ ;
 wire \soc/cpu/cpuregs/_2172_ ;
 wire \soc/cpu/cpuregs/_2173_ ;
 wire \soc/cpu/cpuregs/_2174_ ;
 wire \soc/cpu/cpuregs/_2175_ ;
 wire \soc/cpu/cpuregs/_2176_ ;
 wire \soc/cpu/cpuregs/_2177_ ;
 wire \soc/cpu/cpuregs/_2178_ ;
 wire \soc/cpu/cpuregs/_2179_ ;
 wire \soc/cpu/cpuregs/_2180_ ;
 wire \soc/cpu/cpuregs/_2181_ ;
 wire \soc/cpu/cpuregs/_2182_ ;
 wire \soc/cpu/cpuregs/_2183_ ;
 wire \soc/cpu/cpuregs/_2184_ ;
 wire \soc/cpu/cpuregs/_2185_ ;
 wire \soc/cpu/cpuregs/_2186_ ;
 wire \soc/cpu/cpuregs/_2187_ ;
 wire \soc/cpu/cpuregs/_2188_ ;
 wire \soc/cpu/cpuregs/_2189_ ;
 wire \soc/cpu/cpuregs/_2190_ ;
 wire \soc/cpu/cpuregs/_2191_ ;
 wire \soc/cpu/cpuregs/_2192_ ;
 wire \soc/cpu/cpuregs/_2193_ ;
 wire \soc/cpu/cpuregs/_2194_ ;
 wire \soc/cpu/cpuregs/_2195_ ;
 wire \soc/cpu/cpuregs/_2196_ ;
 wire \soc/cpu/cpuregs/_2197_ ;
 wire \soc/cpu/cpuregs/_2198_ ;
 wire \soc/cpu/cpuregs/_2199_ ;
 wire \soc/cpu/cpuregs/_2200_ ;
 wire \soc/cpu/cpuregs/_2201_ ;
 wire \soc/cpu/cpuregs/_2202_ ;
 wire \soc/cpu/cpuregs/_2203_ ;
 wire \soc/cpu/cpuregs/_2204_ ;
 wire \soc/cpu/cpuregs/_2205_ ;
 wire \soc/cpu/cpuregs/_2206_ ;
 wire \soc/cpu/cpuregs/_2207_ ;
 wire \soc/cpu/cpuregs/_2208_ ;
 wire \soc/cpu/cpuregs/_2209_ ;
 wire \soc/cpu/cpuregs/_2210_ ;
 wire \soc/cpu/cpuregs/_2211_ ;
 wire \soc/cpu/cpuregs/_2212_ ;
 wire \soc/cpu/cpuregs/_2213_ ;
 wire \soc/cpu/cpuregs/_2214_ ;
 wire \soc/cpu/cpuregs/_2215_ ;
 wire \soc/cpu/cpuregs/_2216_ ;
 wire \soc/cpu/cpuregs/_2217_ ;
 wire \soc/cpu/cpuregs/_2218_ ;
 wire \soc/cpu/cpuregs/_2219_ ;
 wire \soc/cpu/cpuregs/_2220_ ;
 wire \soc/cpu/cpuregs/_2221_ ;
 wire \soc/cpu/cpuregs/_2222_ ;
 wire \soc/cpu/cpuregs/_2223_ ;
 wire \soc/cpu/cpuregs/_2224_ ;
 wire \soc/cpu/cpuregs/_2225_ ;
 wire \soc/cpu/cpuregs/_2226_ ;
 wire \soc/cpu/cpuregs/_2227_ ;
 wire \soc/cpu/cpuregs/_2228_ ;
 wire \soc/cpu/cpuregs/_2229_ ;
 wire \soc/cpu/cpuregs/_2230_ ;
 wire \soc/cpu/cpuregs/_2231_ ;
 wire \soc/cpu/cpuregs/_2232_ ;
 wire \soc/cpu/cpuregs/_2233_ ;
 wire \soc/cpu/cpuregs/_2234_ ;
 wire \soc/cpu/cpuregs/_2235_ ;
 wire \soc/cpu/cpuregs/_2236_ ;
 wire \soc/cpu/cpuregs/_2237_ ;
 wire \soc/cpu/cpuregs/_2238_ ;
 wire \soc/cpu/cpuregs/_2239_ ;
 wire \soc/cpu/cpuregs/_2240_ ;
 wire \soc/cpu/cpuregs/_2241_ ;
 wire \soc/cpu/cpuregs/_2242_ ;
 wire \soc/cpu/cpuregs/_2243_ ;
 wire \soc/cpu/cpuregs/_2244_ ;
 wire \soc/cpu/cpuregs/_2245_ ;
 wire \soc/cpu/cpuregs/_2246_ ;
 wire \soc/cpu/cpuregs/_2247_ ;
 wire \soc/cpu/cpuregs/_2248_ ;
 wire \soc/cpu/cpuregs/_2249_ ;
 wire \soc/cpu/cpuregs/_2250_ ;
 wire \soc/cpu/cpuregs/_2251_ ;
 wire \soc/cpu/cpuregs/_2252_ ;
 wire \soc/cpu/cpuregs/_2253_ ;
 wire \soc/cpu/cpuregs/_2254_ ;
 wire \soc/cpu/cpuregs/_2255_ ;
 wire \soc/cpu/cpuregs/_2256_ ;
 wire \soc/cpu/cpuregs/_2257_ ;
 wire \soc/cpu/cpuregs/_2258_ ;
 wire \soc/cpu/cpuregs/_2259_ ;
 wire \soc/cpu/cpuregs/_2260_ ;
 wire \soc/cpu/cpuregs/_2261_ ;
 wire \soc/cpu/cpuregs/_2262_ ;
 wire \soc/cpu/cpuregs/_2263_ ;
 wire \soc/cpu/cpuregs/_2264_ ;
 wire \soc/cpu/cpuregs/_2265_ ;
 wire \soc/cpu/cpuregs/_2266_ ;
 wire \soc/cpu/cpuregs/_2267_ ;
 wire \soc/cpu/cpuregs/_2268_ ;
 wire \soc/cpu/cpuregs/_2269_ ;
 wire \soc/cpu/cpuregs/_2270_ ;
 wire \soc/cpu/cpuregs/_2271_ ;
 wire \soc/cpu/cpuregs/_2272_ ;
 wire \soc/cpu/cpuregs/_2273_ ;
 wire \soc/cpu/cpuregs/_2274_ ;
 wire \soc/cpu/cpuregs/_2275_ ;
 wire clknet_leaf_53_clk;
 wire \soc/cpu/cpuregs/_2277_ ;
 wire \soc/cpu/cpuregs/_2278_ ;
 wire \soc/cpu/cpuregs/_2279_ ;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire \soc/cpu/cpuregs/_2315_ ;
 wire \soc/cpu/cpuregs/_2316_ ;
 wire \soc/cpu/cpuregs/_2317_ ;
 wire \soc/cpu/cpuregs/_2318_ ;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire net491;
 wire net490;
 wire net489;
 wire net487;
 wire net486;
 wire net485;
 wire net484;
 wire net483;
 wire net482;
 wire net481;
 wire net480;
 wire net479;
 wire net478;
 wire net477;
 wire net476;
 wire net475;
 wire net472;
 wire \soc/cpu/cpuregs/_2353_ ;
 wire \soc/cpu/cpuregs/_2354_ ;
 wire \soc/cpu/cpuregs/_2355_ ;
 wire net471;
 wire net470;
 wire net469;
 wire \soc/cpu/cpuregs/_2359_ ;
 wire \soc/cpu/cpuregs/_2360_ ;
 wire \soc/cpu/cpuregs/_2361_ ;
 wire \soc/cpu/cpuregs/_2362_ ;
 wire net468;
 wire net467;
 wire net466;
 wire \soc/cpu/cpuregs/_2366_ ;
 wire \soc/cpu/cpuregs/_2367_ ;
 wire net465;
 wire net464;
 wire net463;
 wire \soc/cpu/cpuregs/_2371_ ;
 wire \soc/cpu/cpuregs/_2372_ ;
 wire \soc/cpu/cpuregs/_2373_ ;
 wire net462;
 wire net461;
 wire net460;
 wire \soc/cpu/cpuregs/_2377_ ;
 wire net459;
 wire net457;
 wire net456;
 wire net455;
 wire \soc/cpu/cpuregs/_2382_ ;
 wire net454;
 wire net453;
 wire net452;
 wire net451;
 wire net450;
 wire net449;
 wire net447;
 wire net446;
 wire net445;
 wire net444;
 wire net443;
 wire net442;
 wire net441;
 wire net440;
 wire net439;
 wire net438;
 wire net437;
 wire net436;
 wire net435;
 wire net434;
 wire net433;
 wire net432;
 wire net431;
 wire net430;
 wire net429;
 wire net428;
 wire net427;
 wire net426;
 wire net425;
 wire net424;
 wire net423;
 wire net422;
 wire net421;
 wire net420;
 wire \soc/cpu/cpuregs/_2417_ ;
 wire net418;
 wire net417;
 wire net416;
 wire \soc/cpu/cpuregs/_2421_ ;
 wire \soc/cpu/cpuregs/_2422_ ;
 wire net415;
 wire net414;
 wire net413;
 wire \soc/cpu/cpuregs/_2426_ ;
 wire \soc/cpu/cpuregs/_2427_ ;
 wire net412;
 wire net411;
 wire net410;
 wire \soc/cpu/cpuregs/_2431_ ;
 wire net409;
 wire net408;
 wire net407;
 wire \soc/cpu/cpuregs/_2435_ ;
 wire \soc/cpu/cpuregs/_2436_ ;
 wire net406;
 wire net405;
 wire net404;
 wire \soc/cpu/cpuregs/_2440_ ;
 wire net403;
 wire net402;
 wire net401;
 wire \soc/cpu/cpuregs/_2444_ ;
 wire net400;
 wire net399;
 wire net398;
 wire \soc/cpu/cpuregs/_2448_ ;
 wire \soc/cpu/cpuregs/_2449_ ;
 wire net397;
 wire net396;
 wire net395;
 wire \soc/cpu/cpuregs/_2453_ ;
 wire \soc/cpu/cpuregs/_2454_ ;
 wire net394;
 wire net393;
 wire net392;
 wire \soc/cpu/cpuregs/_2458_ ;
 wire net391;
 wire net390;
 wire net389;
 wire \soc/cpu/cpuregs/_2462_ ;
 wire net388;
 wire net387;
 wire net386;
 wire \soc/cpu/cpuregs/_2466_ ;
 wire net385;
 wire net384;
 wire net383;
 wire \soc/cpu/cpuregs/_2470_ ;
 wire net382;
 wire net381;
 wire net380;
 wire \soc/cpu/cpuregs/_2474_ ;
 wire net379;
 wire net378;
 wire net377;
 wire \soc/cpu/cpuregs/_2478_ ;
 wire \soc/cpu/cpuregs/_2479_ ;
 wire net376;
 wire net375;
 wire net374;
 wire \soc/cpu/cpuregs/_2483_ ;
 wire net373;
 wire net372;
 wire net371;
 wire \soc/cpu/cpuregs/_2487_ ;
 wire net370;
 wire net369;
 wire net368;
 wire \soc/cpu/cpuregs/_2491_ ;
 wire net367;
 wire net366;
 wire net365;
 wire \soc/cpu/cpuregs/_2495_ ;
 wire net364;
 wire net363;
 wire net362;
 wire \soc/cpu/cpuregs/_2499_ ;
 wire net361;
 wire net360;
 wire net359;
 wire \soc/cpu/cpuregs/_2503_ ;
 wire net358;
 wire net357;
 wire net356;
 wire \soc/cpu/cpuregs/_2507_ ;
 wire net355;
 wire net354;
 wire net353;
 wire \soc/cpu/cpuregs/_2511_ ;
 wire net352;
 wire net351;
 wire net350;
 wire \soc/cpu/cpuregs/_2515_ ;
 wire net349;
 wire net348;
 wire net347;
 wire \soc/cpu/cpuregs/regs[0][0] ;
 wire \soc/cpu/cpuregs/regs[0][10] ;
 wire \soc/cpu/cpuregs/regs[0][11] ;
 wire \soc/cpu/cpuregs/regs[0][12] ;
 wire \soc/cpu/cpuregs/regs[0][13] ;
 wire \soc/cpu/cpuregs/regs[0][14] ;
 wire \soc/cpu/cpuregs/regs[0][15] ;
 wire \soc/cpu/cpuregs/regs[0][16] ;
 wire \soc/cpu/cpuregs/regs[0][17] ;
 wire \soc/cpu/cpuregs/regs[0][18] ;
 wire \soc/cpu/cpuregs/regs[0][19] ;
 wire \soc/cpu/cpuregs/regs[0][1] ;
 wire \soc/cpu/cpuregs/regs[0][20] ;
 wire \soc/cpu/cpuregs/regs[0][21] ;
 wire \soc/cpu/cpuregs/regs[0][22] ;
 wire \soc/cpu/cpuregs/regs[0][23] ;
 wire \soc/cpu/cpuregs/regs[0][24] ;
 wire \soc/cpu/cpuregs/regs[0][25] ;
 wire \soc/cpu/cpuregs/regs[0][26] ;
 wire \soc/cpu/cpuregs/regs[0][27] ;
 wire \soc/cpu/cpuregs/regs[0][28] ;
 wire \soc/cpu/cpuregs/regs[0][29] ;
 wire \soc/cpu/cpuregs/regs[0][2] ;
 wire \soc/cpu/cpuregs/regs[0][30] ;
 wire \soc/cpu/cpuregs/regs[0][31] ;
 wire \soc/cpu/cpuregs/regs[0][3] ;
 wire \soc/cpu/cpuregs/regs[0][4] ;
 wire \soc/cpu/cpuregs/regs[0][5] ;
 wire \soc/cpu/cpuregs/regs[0][6] ;
 wire \soc/cpu/cpuregs/regs[0][7] ;
 wire \soc/cpu/cpuregs/regs[0][8] ;
 wire \soc/cpu/cpuregs/regs[0][9] ;
 wire \soc/cpu/cpuregs/regs[10][0] ;
 wire \soc/cpu/cpuregs/regs[10][10] ;
 wire \soc/cpu/cpuregs/regs[10][11] ;
 wire \soc/cpu/cpuregs/regs[10][12] ;
 wire \soc/cpu/cpuregs/regs[10][13] ;
 wire \soc/cpu/cpuregs/regs[10][14] ;
 wire \soc/cpu/cpuregs/regs[10][15] ;
 wire \soc/cpu/cpuregs/regs[10][16] ;
 wire \soc/cpu/cpuregs/regs[10][17] ;
 wire \soc/cpu/cpuregs/regs[10][18] ;
 wire \soc/cpu/cpuregs/regs[10][19] ;
 wire \soc/cpu/cpuregs/regs[10][1] ;
 wire \soc/cpu/cpuregs/regs[10][20] ;
 wire \soc/cpu/cpuregs/regs[10][21] ;
 wire \soc/cpu/cpuregs/regs[10][22] ;
 wire \soc/cpu/cpuregs/regs[10][23] ;
 wire \soc/cpu/cpuregs/regs[10][24] ;
 wire \soc/cpu/cpuregs/regs[10][25] ;
 wire \soc/cpu/cpuregs/regs[10][26] ;
 wire \soc/cpu/cpuregs/regs[10][27] ;
 wire \soc/cpu/cpuregs/regs[10][28] ;
 wire \soc/cpu/cpuregs/regs[10][29] ;
 wire \soc/cpu/cpuregs/regs[10][2] ;
 wire \soc/cpu/cpuregs/regs[10][30] ;
 wire \soc/cpu/cpuregs/regs[10][31] ;
 wire \soc/cpu/cpuregs/regs[10][3] ;
 wire \soc/cpu/cpuregs/regs[10][4] ;
 wire \soc/cpu/cpuregs/regs[10][5] ;
 wire \soc/cpu/cpuregs/regs[10][6] ;
 wire \soc/cpu/cpuregs/regs[10][7] ;
 wire \soc/cpu/cpuregs/regs[10][8] ;
 wire \soc/cpu/cpuregs/regs[10][9] ;
 wire \soc/cpu/cpuregs/regs[11][0] ;
 wire \soc/cpu/cpuregs/regs[11][10] ;
 wire \soc/cpu/cpuregs/regs[11][11] ;
 wire \soc/cpu/cpuregs/regs[11][12] ;
 wire \soc/cpu/cpuregs/regs[11][13] ;
 wire \soc/cpu/cpuregs/regs[11][14] ;
 wire \soc/cpu/cpuregs/regs[11][15] ;
 wire \soc/cpu/cpuregs/regs[11][16] ;
 wire \soc/cpu/cpuregs/regs[11][17] ;
 wire \soc/cpu/cpuregs/regs[11][18] ;
 wire \soc/cpu/cpuregs/regs[11][19] ;
 wire \soc/cpu/cpuregs/regs[11][1] ;
 wire \soc/cpu/cpuregs/regs[11][20] ;
 wire \soc/cpu/cpuregs/regs[11][21] ;
 wire \soc/cpu/cpuregs/regs[11][22] ;
 wire \soc/cpu/cpuregs/regs[11][23] ;
 wire \soc/cpu/cpuregs/regs[11][24] ;
 wire \soc/cpu/cpuregs/regs[11][25] ;
 wire \soc/cpu/cpuregs/regs[11][26] ;
 wire \soc/cpu/cpuregs/regs[11][27] ;
 wire \soc/cpu/cpuregs/regs[11][28] ;
 wire \soc/cpu/cpuregs/regs[11][29] ;
 wire \soc/cpu/cpuregs/regs[11][2] ;
 wire \soc/cpu/cpuregs/regs[11][30] ;
 wire \soc/cpu/cpuregs/regs[11][31] ;
 wire \soc/cpu/cpuregs/regs[11][3] ;
 wire \soc/cpu/cpuregs/regs[11][4] ;
 wire \soc/cpu/cpuregs/regs[11][5] ;
 wire \soc/cpu/cpuregs/regs[11][6] ;
 wire \soc/cpu/cpuregs/regs[11][7] ;
 wire \soc/cpu/cpuregs/regs[11][8] ;
 wire \soc/cpu/cpuregs/regs[11][9] ;
 wire \soc/cpu/cpuregs/regs[12][0] ;
 wire \soc/cpu/cpuregs/regs[12][10] ;
 wire \soc/cpu/cpuregs/regs[12][11] ;
 wire \soc/cpu/cpuregs/regs[12][12] ;
 wire \soc/cpu/cpuregs/regs[12][13] ;
 wire \soc/cpu/cpuregs/regs[12][14] ;
 wire \soc/cpu/cpuregs/regs[12][15] ;
 wire \soc/cpu/cpuregs/regs[12][16] ;
 wire \soc/cpu/cpuregs/regs[12][17] ;
 wire \soc/cpu/cpuregs/regs[12][18] ;
 wire \soc/cpu/cpuregs/regs[12][19] ;
 wire \soc/cpu/cpuregs/regs[12][1] ;
 wire \soc/cpu/cpuregs/regs[12][20] ;
 wire \soc/cpu/cpuregs/regs[12][21] ;
 wire \soc/cpu/cpuregs/regs[12][22] ;
 wire \soc/cpu/cpuregs/regs[12][23] ;
 wire \soc/cpu/cpuregs/regs[12][24] ;
 wire \soc/cpu/cpuregs/regs[12][25] ;
 wire \soc/cpu/cpuregs/regs[12][26] ;
 wire \soc/cpu/cpuregs/regs[12][27] ;
 wire \soc/cpu/cpuregs/regs[12][28] ;
 wire \soc/cpu/cpuregs/regs[12][29] ;
 wire \soc/cpu/cpuregs/regs[12][2] ;
 wire \soc/cpu/cpuregs/regs[12][30] ;
 wire \soc/cpu/cpuregs/regs[12][31] ;
 wire \soc/cpu/cpuregs/regs[12][3] ;
 wire \soc/cpu/cpuregs/regs[12][4] ;
 wire \soc/cpu/cpuregs/regs[12][5] ;
 wire \soc/cpu/cpuregs/regs[12][6] ;
 wire \soc/cpu/cpuregs/regs[12][7] ;
 wire \soc/cpu/cpuregs/regs[12][8] ;
 wire \soc/cpu/cpuregs/regs[12][9] ;
 wire \soc/cpu/cpuregs/regs[13][0] ;
 wire \soc/cpu/cpuregs/regs[13][10] ;
 wire \soc/cpu/cpuregs/regs[13][11] ;
 wire \soc/cpu/cpuregs/regs[13][12] ;
 wire \soc/cpu/cpuregs/regs[13][13] ;
 wire \soc/cpu/cpuregs/regs[13][14] ;
 wire \soc/cpu/cpuregs/regs[13][15] ;
 wire \soc/cpu/cpuregs/regs[13][16] ;
 wire \soc/cpu/cpuregs/regs[13][17] ;
 wire \soc/cpu/cpuregs/regs[13][18] ;
 wire \soc/cpu/cpuregs/regs[13][19] ;
 wire \soc/cpu/cpuregs/regs[13][1] ;
 wire \soc/cpu/cpuregs/regs[13][20] ;
 wire \soc/cpu/cpuregs/regs[13][21] ;
 wire \soc/cpu/cpuregs/regs[13][22] ;
 wire \soc/cpu/cpuregs/regs[13][23] ;
 wire \soc/cpu/cpuregs/regs[13][24] ;
 wire \soc/cpu/cpuregs/regs[13][25] ;
 wire \soc/cpu/cpuregs/regs[13][26] ;
 wire \soc/cpu/cpuregs/regs[13][27] ;
 wire \soc/cpu/cpuregs/regs[13][28] ;
 wire \soc/cpu/cpuregs/regs[13][29] ;
 wire \soc/cpu/cpuregs/regs[13][2] ;
 wire \soc/cpu/cpuregs/regs[13][30] ;
 wire \soc/cpu/cpuregs/regs[13][31] ;
 wire \soc/cpu/cpuregs/regs[13][3] ;
 wire \soc/cpu/cpuregs/regs[13][4] ;
 wire \soc/cpu/cpuregs/regs[13][5] ;
 wire \soc/cpu/cpuregs/regs[13][6] ;
 wire \soc/cpu/cpuregs/regs[13][7] ;
 wire \soc/cpu/cpuregs/regs[13][8] ;
 wire \soc/cpu/cpuregs/regs[13][9] ;
 wire \soc/cpu/cpuregs/regs[14][0] ;
 wire \soc/cpu/cpuregs/regs[14][10] ;
 wire \soc/cpu/cpuregs/regs[14][11] ;
 wire \soc/cpu/cpuregs/regs[14][12] ;
 wire \soc/cpu/cpuregs/regs[14][13] ;
 wire \soc/cpu/cpuregs/regs[14][14] ;
 wire \soc/cpu/cpuregs/regs[14][15] ;
 wire \soc/cpu/cpuregs/regs[14][16] ;
 wire \soc/cpu/cpuregs/regs[14][17] ;
 wire \soc/cpu/cpuregs/regs[14][18] ;
 wire \soc/cpu/cpuregs/regs[14][19] ;
 wire \soc/cpu/cpuregs/regs[14][1] ;
 wire \soc/cpu/cpuregs/regs[14][20] ;
 wire \soc/cpu/cpuregs/regs[14][21] ;
 wire \soc/cpu/cpuregs/regs[14][22] ;
 wire \soc/cpu/cpuregs/regs[14][23] ;
 wire \soc/cpu/cpuregs/regs[14][24] ;
 wire \soc/cpu/cpuregs/regs[14][25] ;
 wire \soc/cpu/cpuregs/regs[14][26] ;
 wire \soc/cpu/cpuregs/regs[14][27] ;
 wire \soc/cpu/cpuregs/regs[14][28] ;
 wire \soc/cpu/cpuregs/regs[14][29] ;
 wire \soc/cpu/cpuregs/regs[14][2] ;
 wire \soc/cpu/cpuregs/regs[14][30] ;
 wire \soc/cpu/cpuregs/regs[14][31] ;
 wire \soc/cpu/cpuregs/regs[14][3] ;
 wire \soc/cpu/cpuregs/regs[14][4] ;
 wire \soc/cpu/cpuregs/regs[14][5] ;
 wire \soc/cpu/cpuregs/regs[14][6] ;
 wire \soc/cpu/cpuregs/regs[14][7] ;
 wire \soc/cpu/cpuregs/regs[14][8] ;
 wire \soc/cpu/cpuregs/regs[14][9] ;
 wire \soc/cpu/cpuregs/regs[15][0] ;
 wire \soc/cpu/cpuregs/regs[15][10] ;
 wire \soc/cpu/cpuregs/regs[15][11] ;
 wire \soc/cpu/cpuregs/regs[15][12] ;
 wire \soc/cpu/cpuregs/regs[15][13] ;
 wire \soc/cpu/cpuregs/regs[15][14] ;
 wire \soc/cpu/cpuregs/regs[15][15] ;
 wire \soc/cpu/cpuregs/regs[15][16] ;
 wire \soc/cpu/cpuregs/regs[15][17] ;
 wire \soc/cpu/cpuregs/regs[15][18] ;
 wire \soc/cpu/cpuregs/regs[15][19] ;
 wire \soc/cpu/cpuregs/regs[15][1] ;
 wire \soc/cpu/cpuregs/regs[15][20] ;
 wire \soc/cpu/cpuregs/regs[15][21] ;
 wire \soc/cpu/cpuregs/regs[15][22] ;
 wire \soc/cpu/cpuregs/regs[15][23] ;
 wire \soc/cpu/cpuregs/regs[15][24] ;
 wire \soc/cpu/cpuregs/regs[15][25] ;
 wire \soc/cpu/cpuregs/regs[15][26] ;
 wire \soc/cpu/cpuregs/regs[15][27] ;
 wire \soc/cpu/cpuregs/regs[15][28] ;
 wire \soc/cpu/cpuregs/regs[15][29] ;
 wire \soc/cpu/cpuregs/regs[15][2] ;
 wire \soc/cpu/cpuregs/regs[15][30] ;
 wire \soc/cpu/cpuregs/regs[15][31] ;
 wire \soc/cpu/cpuregs/regs[15][3] ;
 wire \soc/cpu/cpuregs/regs[15][4] ;
 wire \soc/cpu/cpuregs/regs[15][5] ;
 wire \soc/cpu/cpuregs/regs[15][6] ;
 wire \soc/cpu/cpuregs/regs[15][7] ;
 wire \soc/cpu/cpuregs/regs[15][8] ;
 wire \soc/cpu/cpuregs/regs[15][9] ;
 wire \soc/cpu/cpuregs/regs[16][0] ;
 wire \soc/cpu/cpuregs/regs[16][10] ;
 wire \soc/cpu/cpuregs/regs[16][11] ;
 wire \soc/cpu/cpuregs/regs[16][12] ;
 wire \soc/cpu/cpuregs/regs[16][13] ;
 wire \soc/cpu/cpuregs/regs[16][14] ;
 wire \soc/cpu/cpuregs/regs[16][15] ;
 wire \soc/cpu/cpuregs/regs[16][16] ;
 wire \soc/cpu/cpuregs/regs[16][17] ;
 wire \soc/cpu/cpuregs/regs[16][18] ;
 wire \soc/cpu/cpuregs/regs[16][19] ;
 wire \soc/cpu/cpuregs/regs[16][1] ;
 wire \soc/cpu/cpuregs/regs[16][20] ;
 wire \soc/cpu/cpuregs/regs[16][21] ;
 wire \soc/cpu/cpuregs/regs[16][22] ;
 wire \soc/cpu/cpuregs/regs[16][23] ;
 wire \soc/cpu/cpuregs/regs[16][24] ;
 wire \soc/cpu/cpuregs/regs[16][25] ;
 wire \soc/cpu/cpuregs/regs[16][26] ;
 wire \soc/cpu/cpuregs/regs[16][27] ;
 wire \soc/cpu/cpuregs/regs[16][28] ;
 wire \soc/cpu/cpuregs/regs[16][29] ;
 wire \soc/cpu/cpuregs/regs[16][2] ;
 wire \soc/cpu/cpuregs/regs[16][30] ;
 wire \soc/cpu/cpuregs/regs[16][31] ;
 wire \soc/cpu/cpuregs/regs[16][3] ;
 wire \soc/cpu/cpuregs/regs[16][4] ;
 wire \soc/cpu/cpuregs/regs[16][5] ;
 wire \soc/cpu/cpuregs/regs[16][6] ;
 wire \soc/cpu/cpuregs/regs[16][7] ;
 wire \soc/cpu/cpuregs/regs[16][8] ;
 wire \soc/cpu/cpuregs/regs[16][9] ;
 wire \soc/cpu/cpuregs/regs[17][0] ;
 wire \soc/cpu/cpuregs/regs[17][10] ;
 wire \soc/cpu/cpuregs/regs[17][11] ;
 wire \soc/cpu/cpuregs/regs[17][12] ;
 wire \soc/cpu/cpuregs/regs[17][13] ;
 wire \soc/cpu/cpuregs/regs[17][14] ;
 wire \soc/cpu/cpuregs/regs[17][15] ;
 wire \soc/cpu/cpuregs/regs[17][16] ;
 wire \soc/cpu/cpuregs/regs[17][17] ;
 wire \soc/cpu/cpuregs/regs[17][18] ;
 wire \soc/cpu/cpuregs/regs[17][19] ;
 wire \soc/cpu/cpuregs/regs[17][1] ;
 wire \soc/cpu/cpuregs/regs[17][20] ;
 wire \soc/cpu/cpuregs/regs[17][21] ;
 wire \soc/cpu/cpuregs/regs[17][22] ;
 wire \soc/cpu/cpuregs/regs[17][23] ;
 wire \soc/cpu/cpuregs/regs[17][24] ;
 wire \soc/cpu/cpuregs/regs[17][25] ;
 wire \soc/cpu/cpuregs/regs[17][26] ;
 wire \soc/cpu/cpuregs/regs[17][27] ;
 wire \soc/cpu/cpuregs/regs[17][28] ;
 wire \soc/cpu/cpuregs/regs[17][29] ;
 wire \soc/cpu/cpuregs/regs[17][2] ;
 wire \soc/cpu/cpuregs/regs[17][30] ;
 wire \soc/cpu/cpuregs/regs[17][31] ;
 wire \soc/cpu/cpuregs/regs[17][3] ;
 wire \soc/cpu/cpuregs/regs[17][4] ;
 wire \soc/cpu/cpuregs/regs[17][5] ;
 wire \soc/cpu/cpuregs/regs[17][6] ;
 wire \soc/cpu/cpuregs/regs[17][7] ;
 wire \soc/cpu/cpuregs/regs[17][8] ;
 wire \soc/cpu/cpuregs/regs[17][9] ;
 wire \soc/cpu/cpuregs/regs[18][0] ;
 wire \soc/cpu/cpuregs/regs[18][10] ;
 wire \soc/cpu/cpuregs/regs[18][11] ;
 wire \soc/cpu/cpuregs/regs[18][12] ;
 wire \soc/cpu/cpuregs/regs[18][13] ;
 wire \soc/cpu/cpuregs/regs[18][14] ;
 wire \soc/cpu/cpuregs/regs[18][15] ;
 wire \soc/cpu/cpuregs/regs[18][16] ;
 wire \soc/cpu/cpuregs/regs[18][17] ;
 wire \soc/cpu/cpuregs/regs[18][18] ;
 wire \soc/cpu/cpuregs/regs[18][19] ;
 wire \soc/cpu/cpuregs/regs[18][1] ;
 wire \soc/cpu/cpuregs/regs[18][20] ;
 wire \soc/cpu/cpuregs/regs[18][21] ;
 wire \soc/cpu/cpuregs/regs[18][22] ;
 wire \soc/cpu/cpuregs/regs[18][23] ;
 wire \soc/cpu/cpuregs/regs[18][24] ;
 wire \soc/cpu/cpuregs/regs[18][25] ;
 wire \soc/cpu/cpuregs/regs[18][26] ;
 wire \soc/cpu/cpuregs/regs[18][27] ;
 wire \soc/cpu/cpuregs/regs[18][28] ;
 wire \soc/cpu/cpuregs/regs[18][29] ;
 wire \soc/cpu/cpuregs/regs[18][2] ;
 wire \soc/cpu/cpuregs/regs[18][30] ;
 wire \soc/cpu/cpuregs/regs[18][31] ;
 wire \soc/cpu/cpuregs/regs[18][3] ;
 wire \soc/cpu/cpuregs/regs[18][4] ;
 wire \soc/cpu/cpuregs/regs[18][5] ;
 wire \soc/cpu/cpuregs/regs[18][6] ;
 wire \soc/cpu/cpuregs/regs[18][7] ;
 wire \soc/cpu/cpuregs/regs[18][8] ;
 wire \soc/cpu/cpuregs/regs[18][9] ;
 wire \soc/cpu/cpuregs/regs[19][0] ;
 wire \soc/cpu/cpuregs/regs[19][10] ;
 wire \soc/cpu/cpuregs/regs[19][11] ;
 wire \soc/cpu/cpuregs/regs[19][12] ;
 wire \soc/cpu/cpuregs/regs[19][13] ;
 wire \soc/cpu/cpuregs/regs[19][14] ;
 wire \soc/cpu/cpuregs/regs[19][15] ;
 wire \soc/cpu/cpuregs/regs[19][16] ;
 wire \soc/cpu/cpuregs/regs[19][17] ;
 wire \soc/cpu/cpuregs/regs[19][18] ;
 wire \soc/cpu/cpuregs/regs[19][19] ;
 wire \soc/cpu/cpuregs/regs[19][1] ;
 wire \soc/cpu/cpuregs/regs[19][20] ;
 wire \soc/cpu/cpuregs/regs[19][21] ;
 wire \soc/cpu/cpuregs/regs[19][22] ;
 wire \soc/cpu/cpuregs/regs[19][23] ;
 wire \soc/cpu/cpuregs/regs[19][24] ;
 wire \soc/cpu/cpuregs/regs[19][25] ;
 wire \soc/cpu/cpuregs/regs[19][26] ;
 wire \soc/cpu/cpuregs/regs[19][27] ;
 wire \soc/cpu/cpuregs/regs[19][28] ;
 wire \soc/cpu/cpuregs/regs[19][29] ;
 wire \soc/cpu/cpuregs/regs[19][2] ;
 wire \soc/cpu/cpuregs/regs[19][30] ;
 wire \soc/cpu/cpuregs/regs[19][31] ;
 wire \soc/cpu/cpuregs/regs[19][3] ;
 wire \soc/cpu/cpuregs/regs[19][4] ;
 wire \soc/cpu/cpuregs/regs[19][5] ;
 wire \soc/cpu/cpuregs/regs[19][6] ;
 wire \soc/cpu/cpuregs/regs[19][7] ;
 wire \soc/cpu/cpuregs/regs[19][8] ;
 wire \soc/cpu/cpuregs/regs[19][9] ;
 wire \soc/cpu/cpuregs/regs[1][0] ;
 wire \soc/cpu/cpuregs/regs[1][10] ;
 wire \soc/cpu/cpuregs/regs[1][11] ;
 wire \soc/cpu/cpuregs/regs[1][12] ;
 wire \soc/cpu/cpuregs/regs[1][13] ;
 wire \soc/cpu/cpuregs/regs[1][14] ;
 wire \soc/cpu/cpuregs/regs[1][15] ;
 wire \soc/cpu/cpuregs/regs[1][16] ;
 wire \soc/cpu/cpuregs/regs[1][17] ;
 wire \soc/cpu/cpuregs/regs[1][18] ;
 wire \soc/cpu/cpuregs/regs[1][19] ;
 wire \soc/cpu/cpuregs/regs[1][1] ;
 wire \soc/cpu/cpuregs/regs[1][20] ;
 wire \soc/cpu/cpuregs/regs[1][21] ;
 wire \soc/cpu/cpuregs/regs[1][22] ;
 wire \soc/cpu/cpuregs/regs[1][23] ;
 wire \soc/cpu/cpuregs/regs[1][24] ;
 wire \soc/cpu/cpuregs/regs[1][25] ;
 wire \soc/cpu/cpuregs/regs[1][26] ;
 wire \soc/cpu/cpuregs/regs[1][27] ;
 wire \soc/cpu/cpuregs/regs[1][28] ;
 wire \soc/cpu/cpuregs/regs[1][29] ;
 wire \soc/cpu/cpuregs/regs[1][2] ;
 wire \soc/cpu/cpuregs/regs[1][30] ;
 wire \soc/cpu/cpuregs/regs[1][31] ;
 wire \soc/cpu/cpuregs/regs[1][3] ;
 wire \soc/cpu/cpuregs/regs[1][4] ;
 wire \soc/cpu/cpuregs/regs[1][5] ;
 wire \soc/cpu/cpuregs/regs[1][6] ;
 wire \soc/cpu/cpuregs/regs[1][7] ;
 wire \soc/cpu/cpuregs/regs[1][8] ;
 wire \soc/cpu/cpuregs/regs[1][9] ;
 wire \soc/cpu/cpuregs/regs[20][0] ;
 wire \soc/cpu/cpuregs/regs[20][10] ;
 wire \soc/cpu/cpuregs/regs[20][11] ;
 wire \soc/cpu/cpuregs/regs[20][12] ;
 wire \soc/cpu/cpuregs/regs[20][13] ;
 wire \soc/cpu/cpuregs/regs[20][14] ;
 wire \soc/cpu/cpuregs/regs[20][15] ;
 wire \soc/cpu/cpuregs/regs[20][16] ;
 wire \soc/cpu/cpuregs/regs[20][17] ;
 wire \soc/cpu/cpuregs/regs[20][18] ;
 wire \soc/cpu/cpuregs/regs[20][19] ;
 wire \soc/cpu/cpuregs/regs[20][1] ;
 wire \soc/cpu/cpuregs/regs[20][20] ;
 wire \soc/cpu/cpuregs/regs[20][21] ;
 wire \soc/cpu/cpuregs/regs[20][22] ;
 wire \soc/cpu/cpuregs/regs[20][23] ;
 wire \soc/cpu/cpuregs/regs[20][24] ;
 wire \soc/cpu/cpuregs/regs[20][25] ;
 wire \soc/cpu/cpuregs/regs[20][26] ;
 wire \soc/cpu/cpuregs/regs[20][27] ;
 wire \soc/cpu/cpuregs/regs[20][28] ;
 wire \soc/cpu/cpuregs/regs[20][29] ;
 wire \soc/cpu/cpuregs/regs[20][2] ;
 wire \soc/cpu/cpuregs/regs[20][30] ;
 wire \soc/cpu/cpuregs/regs[20][31] ;
 wire \soc/cpu/cpuregs/regs[20][3] ;
 wire \soc/cpu/cpuregs/regs[20][4] ;
 wire \soc/cpu/cpuregs/regs[20][5] ;
 wire \soc/cpu/cpuregs/regs[20][6] ;
 wire \soc/cpu/cpuregs/regs[20][7] ;
 wire \soc/cpu/cpuregs/regs[20][8] ;
 wire \soc/cpu/cpuregs/regs[20][9] ;
 wire \soc/cpu/cpuregs/regs[21][0] ;
 wire \soc/cpu/cpuregs/regs[21][10] ;
 wire \soc/cpu/cpuregs/regs[21][11] ;
 wire \soc/cpu/cpuregs/regs[21][12] ;
 wire \soc/cpu/cpuregs/regs[21][13] ;
 wire \soc/cpu/cpuregs/regs[21][14] ;
 wire \soc/cpu/cpuregs/regs[21][15] ;
 wire \soc/cpu/cpuregs/regs[21][16] ;
 wire \soc/cpu/cpuregs/regs[21][17] ;
 wire \soc/cpu/cpuregs/regs[21][18] ;
 wire \soc/cpu/cpuregs/regs[21][19] ;
 wire \soc/cpu/cpuregs/regs[21][1] ;
 wire \soc/cpu/cpuregs/regs[21][20] ;
 wire \soc/cpu/cpuregs/regs[21][21] ;
 wire \soc/cpu/cpuregs/regs[21][22] ;
 wire \soc/cpu/cpuregs/regs[21][23] ;
 wire \soc/cpu/cpuregs/regs[21][24] ;
 wire \soc/cpu/cpuregs/regs[21][25] ;
 wire \soc/cpu/cpuregs/regs[21][26] ;
 wire \soc/cpu/cpuregs/regs[21][27] ;
 wire \soc/cpu/cpuregs/regs[21][28] ;
 wire \soc/cpu/cpuregs/regs[21][29] ;
 wire \soc/cpu/cpuregs/regs[21][2] ;
 wire \soc/cpu/cpuregs/regs[21][30] ;
 wire \soc/cpu/cpuregs/regs[21][31] ;
 wire \soc/cpu/cpuregs/regs[21][3] ;
 wire \soc/cpu/cpuregs/regs[21][4] ;
 wire \soc/cpu/cpuregs/regs[21][5] ;
 wire \soc/cpu/cpuregs/regs[21][6] ;
 wire \soc/cpu/cpuregs/regs[21][7] ;
 wire \soc/cpu/cpuregs/regs[21][8] ;
 wire \soc/cpu/cpuregs/regs[21][9] ;
 wire \soc/cpu/cpuregs/regs[22][0] ;
 wire \soc/cpu/cpuregs/regs[22][10] ;
 wire \soc/cpu/cpuregs/regs[22][11] ;
 wire \soc/cpu/cpuregs/regs[22][12] ;
 wire \soc/cpu/cpuregs/regs[22][13] ;
 wire \soc/cpu/cpuregs/regs[22][14] ;
 wire \soc/cpu/cpuregs/regs[22][15] ;
 wire \soc/cpu/cpuregs/regs[22][16] ;
 wire \soc/cpu/cpuregs/regs[22][17] ;
 wire \soc/cpu/cpuregs/regs[22][18] ;
 wire \soc/cpu/cpuregs/regs[22][19] ;
 wire \soc/cpu/cpuregs/regs[22][1] ;
 wire \soc/cpu/cpuregs/regs[22][20] ;
 wire \soc/cpu/cpuregs/regs[22][21] ;
 wire \soc/cpu/cpuregs/regs[22][22] ;
 wire \soc/cpu/cpuregs/regs[22][23] ;
 wire \soc/cpu/cpuregs/regs[22][24] ;
 wire \soc/cpu/cpuregs/regs[22][25] ;
 wire \soc/cpu/cpuregs/regs[22][26] ;
 wire \soc/cpu/cpuregs/regs[22][27] ;
 wire \soc/cpu/cpuregs/regs[22][28] ;
 wire \soc/cpu/cpuregs/regs[22][29] ;
 wire \soc/cpu/cpuregs/regs[22][2] ;
 wire \soc/cpu/cpuregs/regs[22][30] ;
 wire \soc/cpu/cpuregs/regs[22][31] ;
 wire \soc/cpu/cpuregs/regs[22][3] ;
 wire \soc/cpu/cpuregs/regs[22][4] ;
 wire \soc/cpu/cpuregs/regs[22][5] ;
 wire \soc/cpu/cpuregs/regs[22][6] ;
 wire \soc/cpu/cpuregs/regs[22][7] ;
 wire \soc/cpu/cpuregs/regs[22][8] ;
 wire \soc/cpu/cpuregs/regs[22][9] ;
 wire \soc/cpu/cpuregs/regs[23][0] ;
 wire \soc/cpu/cpuregs/regs[23][10] ;
 wire \soc/cpu/cpuregs/regs[23][11] ;
 wire \soc/cpu/cpuregs/regs[23][12] ;
 wire \soc/cpu/cpuregs/regs[23][13] ;
 wire \soc/cpu/cpuregs/regs[23][14] ;
 wire \soc/cpu/cpuregs/regs[23][15] ;
 wire \soc/cpu/cpuregs/regs[23][16] ;
 wire \soc/cpu/cpuregs/regs[23][17] ;
 wire \soc/cpu/cpuregs/regs[23][18] ;
 wire \soc/cpu/cpuregs/regs[23][19] ;
 wire \soc/cpu/cpuregs/regs[23][1] ;
 wire \soc/cpu/cpuregs/regs[23][20] ;
 wire \soc/cpu/cpuregs/regs[23][21] ;
 wire \soc/cpu/cpuregs/regs[23][22] ;
 wire \soc/cpu/cpuregs/regs[23][23] ;
 wire \soc/cpu/cpuregs/regs[23][24] ;
 wire \soc/cpu/cpuregs/regs[23][25] ;
 wire \soc/cpu/cpuregs/regs[23][26] ;
 wire \soc/cpu/cpuregs/regs[23][27] ;
 wire \soc/cpu/cpuregs/regs[23][28] ;
 wire \soc/cpu/cpuregs/regs[23][29] ;
 wire \soc/cpu/cpuregs/regs[23][2] ;
 wire \soc/cpu/cpuregs/regs[23][30] ;
 wire \soc/cpu/cpuregs/regs[23][31] ;
 wire \soc/cpu/cpuregs/regs[23][3] ;
 wire \soc/cpu/cpuregs/regs[23][4] ;
 wire \soc/cpu/cpuregs/regs[23][5] ;
 wire \soc/cpu/cpuregs/regs[23][6] ;
 wire \soc/cpu/cpuregs/regs[23][7] ;
 wire \soc/cpu/cpuregs/regs[23][8] ;
 wire \soc/cpu/cpuregs/regs[23][9] ;
 wire \soc/cpu/cpuregs/regs[24][0] ;
 wire \soc/cpu/cpuregs/regs[24][10] ;
 wire \soc/cpu/cpuregs/regs[24][11] ;
 wire \soc/cpu/cpuregs/regs[24][12] ;
 wire \soc/cpu/cpuregs/regs[24][13] ;
 wire \soc/cpu/cpuregs/regs[24][14] ;
 wire \soc/cpu/cpuregs/regs[24][15] ;
 wire \soc/cpu/cpuregs/regs[24][16] ;
 wire \soc/cpu/cpuregs/regs[24][17] ;
 wire \soc/cpu/cpuregs/regs[24][18] ;
 wire \soc/cpu/cpuregs/regs[24][19] ;
 wire \soc/cpu/cpuregs/regs[24][1] ;
 wire \soc/cpu/cpuregs/regs[24][20] ;
 wire \soc/cpu/cpuregs/regs[24][21] ;
 wire \soc/cpu/cpuregs/regs[24][22] ;
 wire \soc/cpu/cpuregs/regs[24][23] ;
 wire \soc/cpu/cpuregs/regs[24][24] ;
 wire \soc/cpu/cpuregs/regs[24][25] ;
 wire \soc/cpu/cpuregs/regs[24][26] ;
 wire \soc/cpu/cpuregs/regs[24][27] ;
 wire \soc/cpu/cpuregs/regs[24][28] ;
 wire \soc/cpu/cpuregs/regs[24][29] ;
 wire \soc/cpu/cpuregs/regs[24][2] ;
 wire \soc/cpu/cpuregs/regs[24][30] ;
 wire \soc/cpu/cpuregs/regs[24][31] ;
 wire \soc/cpu/cpuregs/regs[24][3] ;
 wire \soc/cpu/cpuregs/regs[24][4] ;
 wire \soc/cpu/cpuregs/regs[24][5] ;
 wire \soc/cpu/cpuregs/regs[24][6] ;
 wire \soc/cpu/cpuregs/regs[24][7] ;
 wire \soc/cpu/cpuregs/regs[24][8] ;
 wire \soc/cpu/cpuregs/regs[24][9] ;
 wire \soc/cpu/cpuregs/regs[25][0] ;
 wire \soc/cpu/cpuregs/regs[25][10] ;
 wire \soc/cpu/cpuregs/regs[25][11] ;
 wire \soc/cpu/cpuregs/regs[25][12] ;
 wire \soc/cpu/cpuregs/regs[25][13] ;
 wire \soc/cpu/cpuregs/regs[25][14] ;
 wire \soc/cpu/cpuregs/regs[25][15] ;
 wire \soc/cpu/cpuregs/regs[25][16] ;
 wire \soc/cpu/cpuregs/regs[25][17] ;
 wire \soc/cpu/cpuregs/regs[25][18] ;
 wire \soc/cpu/cpuregs/regs[25][19] ;
 wire \soc/cpu/cpuregs/regs[25][1] ;
 wire \soc/cpu/cpuregs/regs[25][20] ;
 wire \soc/cpu/cpuregs/regs[25][21] ;
 wire \soc/cpu/cpuregs/regs[25][22] ;
 wire \soc/cpu/cpuregs/regs[25][23] ;
 wire \soc/cpu/cpuregs/regs[25][24] ;
 wire \soc/cpu/cpuregs/regs[25][25] ;
 wire \soc/cpu/cpuregs/regs[25][26] ;
 wire \soc/cpu/cpuregs/regs[25][27] ;
 wire \soc/cpu/cpuregs/regs[25][28] ;
 wire \soc/cpu/cpuregs/regs[25][29] ;
 wire \soc/cpu/cpuregs/regs[25][2] ;
 wire \soc/cpu/cpuregs/regs[25][30] ;
 wire \soc/cpu/cpuregs/regs[25][31] ;
 wire \soc/cpu/cpuregs/regs[25][3] ;
 wire \soc/cpu/cpuregs/regs[25][4] ;
 wire \soc/cpu/cpuregs/regs[25][5] ;
 wire \soc/cpu/cpuregs/regs[25][6] ;
 wire \soc/cpu/cpuregs/regs[25][7] ;
 wire \soc/cpu/cpuregs/regs[25][8] ;
 wire \soc/cpu/cpuregs/regs[25][9] ;
 wire \soc/cpu/cpuregs/regs[26][0] ;
 wire \soc/cpu/cpuregs/regs[26][10] ;
 wire \soc/cpu/cpuregs/regs[26][11] ;
 wire \soc/cpu/cpuregs/regs[26][12] ;
 wire \soc/cpu/cpuregs/regs[26][13] ;
 wire \soc/cpu/cpuregs/regs[26][14] ;
 wire \soc/cpu/cpuregs/regs[26][15] ;
 wire \soc/cpu/cpuregs/regs[26][16] ;
 wire \soc/cpu/cpuregs/regs[26][17] ;
 wire \soc/cpu/cpuregs/regs[26][18] ;
 wire \soc/cpu/cpuregs/regs[26][19] ;
 wire \soc/cpu/cpuregs/regs[26][1] ;
 wire \soc/cpu/cpuregs/regs[26][20] ;
 wire \soc/cpu/cpuregs/regs[26][21] ;
 wire \soc/cpu/cpuregs/regs[26][22] ;
 wire \soc/cpu/cpuregs/regs[26][23] ;
 wire \soc/cpu/cpuregs/regs[26][24] ;
 wire \soc/cpu/cpuregs/regs[26][25] ;
 wire \soc/cpu/cpuregs/regs[26][26] ;
 wire \soc/cpu/cpuregs/regs[26][27] ;
 wire \soc/cpu/cpuregs/regs[26][28] ;
 wire \soc/cpu/cpuregs/regs[26][29] ;
 wire \soc/cpu/cpuregs/regs[26][2] ;
 wire \soc/cpu/cpuregs/regs[26][30] ;
 wire \soc/cpu/cpuregs/regs[26][31] ;
 wire \soc/cpu/cpuregs/regs[26][3] ;
 wire \soc/cpu/cpuregs/regs[26][4] ;
 wire \soc/cpu/cpuregs/regs[26][5] ;
 wire \soc/cpu/cpuregs/regs[26][6] ;
 wire \soc/cpu/cpuregs/regs[26][7] ;
 wire \soc/cpu/cpuregs/regs[26][8] ;
 wire \soc/cpu/cpuregs/regs[26][9] ;
 wire \soc/cpu/cpuregs/regs[27][0] ;
 wire \soc/cpu/cpuregs/regs[27][10] ;
 wire \soc/cpu/cpuregs/regs[27][11] ;
 wire \soc/cpu/cpuregs/regs[27][12] ;
 wire \soc/cpu/cpuregs/regs[27][13] ;
 wire \soc/cpu/cpuregs/regs[27][14] ;
 wire \soc/cpu/cpuregs/regs[27][15] ;
 wire \soc/cpu/cpuregs/regs[27][16] ;
 wire \soc/cpu/cpuregs/regs[27][17] ;
 wire \soc/cpu/cpuregs/regs[27][18] ;
 wire \soc/cpu/cpuregs/regs[27][19] ;
 wire \soc/cpu/cpuregs/regs[27][1] ;
 wire \soc/cpu/cpuregs/regs[27][20] ;
 wire \soc/cpu/cpuregs/regs[27][21] ;
 wire \soc/cpu/cpuregs/regs[27][22] ;
 wire \soc/cpu/cpuregs/regs[27][23] ;
 wire \soc/cpu/cpuregs/regs[27][24] ;
 wire \soc/cpu/cpuregs/regs[27][25] ;
 wire \soc/cpu/cpuregs/regs[27][26] ;
 wire \soc/cpu/cpuregs/regs[27][27] ;
 wire \soc/cpu/cpuregs/regs[27][28] ;
 wire \soc/cpu/cpuregs/regs[27][29] ;
 wire \soc/cpu/cpuregs/regs[27][2] ;
 wire \soc/cpu/cpuregs/regs[27][30] ;
 wire \soc/cpu/cpuregs/regs[27][31] ;
 wire \soc/cpu/cpuregs/regs[27][3] ;
 wire \soc/cpu/cpuregs/regs[27][4] ;
 wire \soc/cpu/cpuregs/regs[27][5] ;
 wire \soc/cpu/cpuregs/regs[27][6] ;
 wire \soc/cpu/cpuregs/regs[27][7] ;
 wire \soc/cpu/cpuregs/regs[27][8] ;
 wire \soc/cpu/cpuregs/regs[27][9] ;
 wire \soc/cpu/cpuregs/regs[28][0] ;
 wire \soc/cpu/cpuregs/regs[28][10] ;
 wire \soc/cpu/cpuregs/regs[28][11] ;
 wire \soc/cpu/cpuregs/regs[28][12] ;
 wire \soc/cpu/cpuregs/regs[28][13] ;
 wire \soc/cpu/cpuregs/regs[28][14] ;
 wire \soc/cpu/cpuregs/regs[28][15] ;
 wire \soc/cpu/cpuregs/regs[28][16] ;
 wire \soc/cpu/cpuregs/regs[28][17] ;
 wire \soc/cpu/cpuregs/regs[28][18] ;
 wire \soc/cpu/cpuregs/regs[28][19] ;
 wire \soc/cpu/cpuregs/regs[28][1] ;
 wire \soc/cpu/cpuregs/regs[28][20] ;
 wire \soc/cpu/cpuregs/regs[28][21] ;
 wire \soc/cpu/cpuregs/regs[28][22] ;
 wire \soc/cpu/cpuregs/regs[28][23] ;
 wire \soc/cpu/cpuregs/regs[28][24] ;
 wire \soc/cpu/cpuregs/regs[28][25] ;
 wire \soc/cpu/cpuregs/regs[28][26] ;
 wire \soc/cpu/cpuregs/regs[28][27] ;
 wire \soc/cpu/cpuregs/regs[28][28] ;
 wire \soc/cpu/cpuregs/regs[28][29] ;
 wire \soc/cpu/cpuregs/regs[28][2] ;
 wire \soc/cpu/cpuregs/regs[28][30] ;
 wire \soc/cpu/cpuregs/regs[28][31] ;
 wire \soc/cpu/cpuregs/regs[28][3] ;
 wire \soc/cpu/cpuregs/regs[28][4] ;
 wire \soc/cpu/cpuregs/regs[28][5] ;
 wire \soc/cpu/cpuregs/regs[28][6] ;
 wire \soc/cpu/cpuregs/regs[28][7] ;
 wire \soc/cpu/cpuregs/regs[28][8] ;
 wire \soc/cpu/cpuregs/regs[28][9] ;
 wire \soc/cpu/cpuregs/regs[29][0] ;
 wire \soc/cpu/cpuregs/regs[29][10] ;
 wire \soc/cpu/cpuregs/regs[29][11] ;
 wire \soc/cpu/cpuregs/regs[29][12] ;
 wire \soc/cpu/cpuregs/regs[29][13] ;
 wire \soc/cpu/cpuregs/regs[29][14] ;
 wire \soc/cpu/cpuregs/regs[29][15] ;
 wire \soc/cpu/cpuregs/regs[29][16] ;
 wire \soc/cpu/cpuregs/regs[29][17] ;
 wire \soc/cpu/cpuregs/regs[29][18] ;
 wire \soc/cpu/cpuregs/regs[29][19] ;
 wire \soc/cpu/cpuregs/regs[29][1] ;
 wire \soc/cpu/cpuregs/regs[29][20] ;
 wire \soc/cpu/cpuregs/regs[29][21] ;
 wire \soc/cpu/cpuregs/regs[29][22] ;
 wire \soc/cpu/cpuregs/regs[29][23] ;
 wire \soc/cpu/cpuregs/regs[29][24] ;
 wire \soc/cpu/cpuregs/regs[29][25] ;
 wire \soc/cpu/cpuregs/regs[29][26] ;
 wire \soc/cpu/cpuregs/regs[29][27] ;
 wire \soc/cpu/cpuregs/regs[29][28] ;
 wire \soc/cpu/cpuregs/regs[29][29] ;
 wire \soc/cpu/cpuregs/regs[29][2] ;
 wire \soc/cpu/cpuregs/regs[29][30] ;
 wire \soc/cpu/cpuregs/regs[29][31] ;
 wire \soc/cpu/cpuregs/regs[29][3] ;
 wire \soc/cpu/cpuregs/regs[29][4] ;
 wire \soc/cpu/cpuregs/regs[29][5] ;
 wire \soc/cpu/cpuregs/regs[29][6] ;
 wire \soc/cpu/cpuregs/regs[29][7] ;
 wire \soc/cpu/cpuregs/regs[29][8] ;
 wire \soc/cpu/cpuregs/regs[29][9] ;
 wire \soc/cpu/cpuregs/regs[2][0] ;
 wire \soc/cpu/cpuregs/regs[2][10] ;
 wire \soc/cpu/cpuregs/regs[2][11] ;
 wire \soc/cpu/cpuregs/regs[2][12] ;
 wire \soc/cpu/cpuregs/regs[2][13] ;
 wire \soc/cpu/cpuregs/regs[2][14] ;
 wire \soc/cpu/cpuregs/regs[2][15] ;
 wire \soc/cpu/cpuregs/regs[2][16] ;
 wire \soc/cpu/cpuregs/regs[2][17] ;
 wire \soc/cpu/cpuregs/regs[2][18] ;
 wire \soc/cpu/cpuregs/regs[2][19] ;
 wire \soc/cpu/cpuregs/regs[2][1] ;
 wire \soc/cpu/cpuregs/regs[2][20] ;
 wire \soc/cpu/cpuregs/regs[2][21] ;
 wire \soc/cpu/cpuregs/regs[2][22] ;
 wire \soc/cpu/cpuregs/regs[2][23] ;
 wire \soc/cpu/cpuregs/regs[2][24] ;
 wire \soc/cpu/cpuregs/regs[2][25] ;
 wire \soc/cpu/cpuregs/regs[2][26] ;
 wire \soc/cpu/cpuregs/regs[2][27] ;
 wire \soc/cpu/cpuregs/regs[2][28] ;
 wire \soc/cpu/cpuregs/regs[2][29] ;
 wire \soc/cpu/cpuregs/regs[2][2] ;
 wire \soc/cpu/cpuregs/regs[2][30] ;
 wire \soc/cpu/cpuregs/regs[2][31] ;
 wire \soc/cpu/cpuregs/regs[2][3] ;
 wire \soc/cpu/cpuregs/regs[2][4] ;
 wire \soc/cpu/cpuregs/regs[2][5] ;
 wire \soc/cpu/cpuregs/regs[2][6] ;
 wire \soc/cpu/cpuregs/regs[2][7] ;
 wire \soc/cpu/cpuregs/regs[2][8] ;
 wire \soc/cpu/cpuregs/regs[2][9] ;
 wire \soc/cpu/cpuregs/regs[30][0] ;
 wire \soc/cpu/cpuregs/regs[30][10] ;
 wire \soc/cpu/cpuregs/regs[30][11] ;
 wire \soc/cpu/cpuregs/regs[30][12] ;
 wire \soc/cpu/cpuregs/regs[30][13] ;
 wire \soc/cpu/cpuregs/regs[30][14] ;
 wire \soc/cpu/cpuregs/regs[30][15] ;
 wire \soc/cpu/cpuregs/regs[30][16] ;
 wire \soc/cpu/cpuregs/regs[30][17] ;
 wire \soc/cpu/cpuregs/regs[30][18] ;
 wire \soc/cpu/cpuregs/regs[30][19] ;
 wire \soc/cpu/cpuregs/regs[30][1] ;
 wire \soc/cpu/cpuregs/regs[30][20] ;
 wire \soc/cpu/cpuregs/regs[30][21] ;
 wire \soc/cpu/cpuregs/regs[30][22] ;
 wire \soc/cpu/cpuregs/regs[30][23] ;
 wire \soc/cpu/cpuregs/regs[30][24] ;
 wire \soc/cpu/cpuregs/regs[30][25] ;
 wire \soc/cpu/cpuregs/regs[30][26] ;
 wire \soc/cpu/cpuregs/regs[30][27] ;
 wire \soc/cpu/cpuregs/regs[30][28] ;
 wire \soc/cpu/cpuregs/regs[30][29] ;
 wire \soc/cpu/cpuregs/regs[30][2] ;
 wire \soc/cpu/cpuregs/regs[30][30] ;
 wire \soc/cpu/cpuregs/regs[30][31] ;
 wire \soc/cpu/cpuregs/regs[30][3] ;
 wire \soc/cpu/cpuregs/regs[30][4] ;
 wire \soc/cpu/cpuregs/regs[30][5] ;
 wire \soc/cpu/cpuregs/regs[30][6] ;
 wire \soc/cpu/cpuregs/regs[30][7] ;
 wire \soc/cpu/cpuregs/regs[30][8] ;
 wire \soc/cpu/cpuregs/regs[30][9] ;
 wire \soc/cpu/cpuregs/regs[31][0] ;
 wire \soc/cpu/cpuregs/regs[31][10] ;
 wire \soc/cpu/cpuregs/regs[31][11] ;
 wire \soc/cpu/cpuregs/regs[31][12] ;
 wire \soc/cpu/cpuregs/regs[31][13] ;
 wire \soc/cpu/cpuregs/regs[31][14] ;
 wire \soc/cpu/cpuregs/regs[31][15] ;
 wire \soc/cpu/cpuregs/regs[31][16] ;
 wire \soc/cpu/cpuregs/regs[31][17] ;
 wire \soc/cpu/cpuregs/regs[31][18] ;
 wire \soc/cpu/cpuregs/regs[31][19] ;
 wire \soc/cpu/cpuregs/regs[31][1] ;
 wire \soc/cpu/cpuregs/regs[31][20] ;
 wire \soc/cpu/cpuregs/regs[31][21] ;
 wire \soc/cpu/cpuregs/regs[31][22] ;
 wire \soc/cpu/cpuregs/regs[31][23] ;
 wire \soc/cpu/cpuregs/regs[31][24] ;
 wire \soc/cpu/cpuregs/regs[31][25] ;
 wire \soc/cpu/cpuregs/regs[31][26] ;
 wire \soc/cpu/cpuregs/regs[31][27] ;
 wire \soc/cpu/cpuregs/regs[31][28] ;
 wire \soc/cpu/cpuregs/regs[31][29] ;
 wire \soc/cpu/cpuregs/regs[31][2] ;
 wire \soc/cpu/cpuregs/regs[31][30] ;
 wire \soc/cpu/cpuregs/regs[31][31] ;
 wire \soc/cpu/cpuregs/regs[31][3] ;
 wire \soc/cpu/cpuregs/regs[31][4] ;
 wire \soc/cpu/cpuregs/regs[31][5] ;
 wire \soc/cpu/cpuregs/regs[31][6] ;
 wire \soc/cpu/cpuregs/regs[31][7] ;
 wire \soc/cpu/cpuregs/regs[31][8] ;
 wire \soc/cpu/cpuregs/regs[31][9] ;
 wire \soc/cpu/cpuregs/regs[3][0] ;
 wire \soc/cpu/cpuregs/regs[3][10] ;
 wire \soc/cpu/cpuregs/regs[3][11] ;
 wire \soc/cpu/cpuregs/regs[3][12] ;
 wire \soc/cpu/cpuregs/regs[3][13] ;
 wire \soc/cpu/cpuregs/regs[3][14] ;
 wire \soc/cpu/cpuregs/regs[3][15] ;
 wire \soc/cpu/cpuregs/regs[3][16] ;
 wire \soc/cpu/cpuregs/regs[3][17] ;
 wire \soc/cpu/cpuregs/regs[3][18] ;
 wire \soc/cpu/cpuregs/regs[3][19] ;
 wire \soc/cpu/cpuregs/regs[3][1] ;
 wire \soc/cpu/cpuregs/regs[3][20] ;
 wire \soc/cpu/cpuregs/regs[3][21] ;
 wire \soc/cpu/cpuregs/regs[3][22] ;
 wire \soc/cpu/cpuregs/regs[3][23] ;
 wire \soc/cpu/cpuregs/regs[3][24] ;
 wire \soc/cpu/cpuregs/regs[3][25] ;
 wire \soc/cpu/cpuregs/regs[3][26] ;
 wire \soc/cpu/cpuregs/regs[3][27] ;
 wire \soc/cpu/cpuregs/regs[3][28] ;
 wire \soc/cpu/cpuregs/regs[3][29] ;
 wire \soc/cpu/cpuregs/regs[3][2] ;
 wire \soc/cpu/cpuregs/regs[3][30] ;
 wire \soc/cpu/cpuregs/regs[3][31] ;
 wire \soc/cpu/cpuregs/regs[3][3] ;
 wire \soc/cpu/cpuregs/regs[3][4] ;
 wire \soc/cpu/cpuregs/regs[3][5] ;
 wire \soc/cpu/cpuregs/regs[3][6] ;
 wire \soc/cpu/cpuregs/regs[3][7] ;
 wire \soc/cpu/cpuregs/regs[3][8] ;
 wire \soc/cpu/cpuregs/regs[3][9] ;
 wire \soc/cpu/cpuregs/regs[4][0] ;
 wire \soc/cpu/cpuregs/regs[4][10] ;
 wire \soc/cpu/cpuregs/regs[4][11] ;
 wire \soc/cpu/cpuregs/regs[4][12] ;
 wire \soc/cpu/cpuregs/regs[4][13] ;
 wire \soc/cpu/cpuregs/regs[4][14] ;
 wire \soc/cpu/cpuregs/regs[4][15] ;
 wire \soc/cpu/cpuregs/regs[4][16] ;
 wire \soc/cpu/cpuregs/regs[4][17] ;
 wire \soc/cpu/cpuregs/regs[4][18] ;
 wire \soc/cpu/cpuregs/regs[4][19] ;
 wire \soc/cpu/cpuregs/regs[4][1] ;
 wire \soc/cpu/cpuregs/regs[4][20] ;
 wire \soc/cpu/cpuregs/regs[4][21] ;
 wire \soc/cpu/cpuregs/regs[4][22] ;
 wire \soc/cpu/cpuregs/regs[4][23] ;
 wire \soc/cpu/cpuregs/regs[4][24] ;
 wire \soc/cpu/cpuregs/regs[4][25] ;
 wire \soc/cpu/cpuregs/regs[4][26] ;
 wire \soc/cpu/cpuregs/regs[4][27] ;
 wire \soc/cpu/cpuregs/regs[4][28] ;
 wire \soc/cpu/cpuregs/regs[4][29] ;
 wire \soc/cpu/cpuregs/regs[4][2] ;
 wire \soc/cpu/cpuregs/regs[4][30] ;
 wire \soc/cpu/cpuregs/regs[4][31] ;
 wire \soc/cpu/cpuregs/regs[4][3] ;
 wire \soc/cpu/cpuregs/regs[4][4] ;
 wire \soc/cpu/cpuregs/regs[4][5] ;
 wire \soc/cpu/cpuregs/regs[4][6] ;
 wire \soc/cpu/cpuregs/regs[4][7] ;
 wire \soc/cpu/cpuregs/regs[4][8] ;
 wire \soc/cpu/cpuregs/regs[4][9] ;
 wire \soc/cpu/cpuregs/regs[5][0] ;
 wire \soc/cpu/cpuregs/regs[5][10] ;
 wire \soc/cpu/cpuregs/regs[5][11] ;
 wire \soc/cpu/cpuregs/regs[5][12] ;
 wire \soc/cpu/cpuregs/regs[5][13] ;
 wire \soc/cpu/cpuregs/regs[5][14] ;
 wire \soc/cpu/cpuregs/regs[5][15] ;
 wire \soc/cpu/cpuregs/regs[5][16] ;
 wire \soc/cpu/cpuregs/regs[5][17] ;
 wire \soc/cpu/cpuregs/regs[5][18] ;
 wire \soc/cpu/cpuregs/regs[5][19] ;
 wire \soc/cpu/cpuregs/regs[5][1] ;
 wire \soc/cpu/cpuregs/regs[5][20] ;
 wire \soc/cpu/cpuregs/regs[5][21] ;
 wire \soc/cpu/cpuregs/regs[5][22] ;
 wire \soc/cpu/cpuregs/regs[5][23] ;
 wire \soc/cpu/cpuregs/regs[5][24] ;
 wire \soc/cpu/cpuregs/regs[5][25] ;
 wire \soc/cpu/cpuregs/regs[5][26] ;
 wire \soc/cpu/cpuregs/regs[5][27] ;
 wire \soc/cpu/cpuregs/regs[5][28] ;
 wire \soc/cpu/cpuregs/regs[5][29] ;
 wire \soc/cpu/cpuregs/regs[5][2] ;
 wire \soc/cpu/cpuregs/regs[5][30] ;
 wire \soc/cpu/cpuregs/regs[5][31] ;
 wire \soc/cpu/cpuregs/regs[5][3] ;
 wire \soc/cpu/cpuregs/regs[5][4] ;
 wire \soc/cpu/cpuregs/regs[5][5] ;
 wire \soc/cpu/cpuregs/regs[5][6] ;
 wire \soc/cpu/cpuregs/regs[5][7] ;
 wire \soc/cpu/cpuregs/regs[5][8] ;
 wire \soc/cpu/cpuregs/regs[5][9] ;
 wire \soc/cpu/cpuregs/regs[6][0] ;
 wire \soc/cpu/cpuregs/regs[6][10] ;
 wire \soc/cpu/cpuregs/regs[6][11] ;
 wire \soc/cpu/cpuregs/regs[6][12] ;
 wire \soc/cpu/cpuregs/regs[6][13] ;
 wire \soc/cpu/cpuregs/regs[6][14] ;
 wire \soc/cpu/cpuregs/regs[6][15] ;
 wire \soc/cpu/cpuregs/regs[6][16] ;
 wire \soc/cpu/cpuregs/regs[6][17] ;
 wire \soc/cpu/cpuregs/regs[6][18] ;
 wire \soc/cpu/cpuregs/regs[6][19] ;
 wire \soc/cpu/cpuregs/regs[6][1] ;
 wire \soc/cpu/cpuregs/regs[6][20] ;
 wire \soc/cpu/cpuregs/regs[6][21] ;
 wire \soc/cpu/cpuregs/regs[6][22] ;
 wire \soc/cpu/cpuregs/regs[6][23] ;
 wire \soc/cpu/cpuregs/regs[6][24] ;
 wire \soc/cpu/cpuregs/regs[6][25] ;
 wire \soc/cpu/cpuregs/regs[6][26] ;
 wire \soc/cpu/cpuregs/regs[6][27] ;
 wire \soc/cpu/cpuregs/regs[6][28] ;
 wire \soc/cpu/cpuregs/regs[6][29] ;
 wire \soc/cpu/cpuregs/regs[6][2] ;
 wire \soc/cpu/cpuregs/regs[6][30] ;
 wire \soc/cpu/cpuregs/regs[6][31] ;
 wire \soc/cpu/cpuregs/regs[6][3] ;
 wire \soc/cpu/cpuregs/regs[6][4] ;
 wire \soc/cpu/cpuregs/regs[6][5] ;
 wire \soc/cpu/cpuregs/regs[6][6] ;
 wire \soc/cpu/cpuregs/regs[6][7] ;
 wire \soc/cpu/cpuregs/regs[6][8] ;
 wire \soc/cpu/cpuregs/regs[6][9] ;
 wire \soc/cpu/cpuregs/regs[7][0] ;
 wire \soc/cpu/cpuregs/regs[7][10] ;
 wire \soc/cpu/cpuregs/regs[7][11] ;
 wire \soc/cpu/cpuregs/regs[7][12] ;
 wire \soc/cpu/cpuregs/regs[7][13] ;
 wire \soc/cpu/cpuregs/regs[7][14] ;
 wire \soc/cpu/cpuregs/regs[7][15] ;
 wire \soc/cpu/cpuregs/regs[7][16] ;
 wire \soc/cpu/cpuregs/regs[7][17] ;
 wire \soc/cpu/cpuregs/regs[7][18] ;
 wire \soc/cpu/cpuregs/regs[7][19] ;
 wire \soc/cpu/cpuregs/regs[7][1] ;
 wire \soc/cpu/cpuregs/regs[7][20] ;
 wire \soc/cpu/cpuregs/regs[7][21] ;
 wire \soc/cpu/cpuregs/regs[7][22] ;
 wire \soc/cpu/cpuregs/regs[7][23] ;
 wire \soc/cpu/cpuregs/regs[7][24] ;
 wire \soc/cpu/cpuregs/regs[7][25] ;
 wire \soc/cpu/cpuregs/regs[7][26] ;
 wire \soc/cpu/cpuregs/regs[7][27] ;
 wire \soc/cpu/cpuregs/regs[7][28] ;
 wire \soc/cpu/cpuregs/regs[7][29] ;
 wire \soc/cpu/cpuregs/regs[7][2] ;
 wire \soc/cpu/cpuregs/regs[7][30] ;
 wire \soc/cpu/cpuregs/regs[7][31] ;
 wire \soc/cpu/cpuregs/regs[7][3] ;
 wire \soc/cpu/cpuregs/regs[7][4] ;
 wire \soc/cpu/cpuregs/regs[7][5] ;
 wire \soc/cpu/cpuregs/regs[7][6] ;
 wire \soc/cpu/cpuregs/regs[7][7] ;
 wire \soc/cpu/cpuregs/regs[7][8] ;
 wire \soc/cpu/cpuregs/regs[7][9] ;
 wire \soc/cpu/cpuregs/regs[8][0] ;
 wire \soc/cpu/cpuregs/regs[8][10] ;
 wire \soc/cpu/cpuregs/regs[8][11] ;
 wire \soc/cpu/cpuregs/regs[8][12] ;
 wire \soc/cpu/cpuregs/regs[8][13] ;
 wire \soc/cpu/cpuregs/regs[8][14] ;
 wire \soc/cpu/cpuregs/regs[8][15] ;
 wire \soc/cpu/cpuregs/regs[8][16] ;
 wire \soc/cpu/cpuregs/regs[8][17] ;
 wire \soc/cpu/cpuregs/regs[8][18] ;
 wire \soc/cpu/cpuregs/regs[8][19] ;
 wire \soc/cpu/cpuregs/regs[8][1] ;
 wire \soc/cpu/cpuregs/regs[8][20] ;
 wire \soc/cpu/cpuregs/regs[8][21] ;
 wire \soc/cpu/cpuregs/regs[8][22] ;
 wire \soc/cpu/cpuregs/regs[8][23] ;
 wire \soc/cpu/cpuregs/regs[8][24] ;
 wire \soc/cpu/cpuregs/regs[8][25] ;
 wire \soc/cpu/cpuregs/regs[8][26] ;
 wire \soc/cpu/cpuregs/regs[8][27] ;
 wire \soc/cpu/cpuregs/regs[8][28] ;
 wire \soc/cpu/cpuregs/regs[8][29] ;
 wire \soc/cpu/cpuregs/regs[8][2] ;
 wire \soc/cpu/cpuregs/regs[8][30] ;
 wire \soc/cpu/cpuregs/regs[8][31] ;
 wire \soc/cpu/cpuregs/regs[8][3] ;
 wire \soc/cpu/cpuregs/regs[8][4] ;
 wire \soc/cpu/cpuregs/regs[8][5] ;
 wire \soc/cpu/cpuregs/regs[8][6] ;
 wire \soc/cpu/cpuregs/regs[8][7] ;
 wire \soc/cpu/cpuregs/regs[8][8] ;
 wire \soc/cpu/cpuregs/regs[8][9] ;
 wire \soc/cpu/cpuregs/regs[9][0] ;
 wire \soc/cpu/cpuregs/regs[9][10] ;
 wire \soc/cpu/cpuregs/regs[9][11] ;
 wire \soc/cpu/cpuregs/regs[9][12] ;
 wire \soc/cpu/cpuregs/regs[9][13] ;
 wire \soc/cpu/cpuregs/regs[9][14] ;
 wire \soc/cpu/cpuregs/regs[9][15] ;
 wire \soc/cpu/cpuregs/regs[9][16] ;
 wire \soc/cpu/cpuregs/regs[9][17] ;
 wire \soc/cpu/cpuregs/regs[9][18] ;
 wire \soc/cpu/cpuregs/regs[9][19] ;
 wire \soc/cpu/cpuregs/regs[9][1] ;
 wire \soc/cpu/cpuregs/regs[9][20] ;
 wire \soc/cpu/cpuregs/regs[9][21] ;
 wire \soc/cpu/cpuregs/regs[9][22] ;
 wire \soc/cpu/cpuregs/regs[9][23] ;
 wire \soc/cpu/cpuregs/regs[9][24] ;
 wire \soc/cpu/cpuregs/regs[9][25] ;
 wire \soc/cpu/cpuregs/regs[9][26] ;
 wire \soc/cpu/cpuregs/regs[9][27] ;
 wire \soc/cpu/cpuregs/regs[9][28] ;
 wire \soc/cpu/cpuregs/regs[9][29] ;
 wire \soc/cpu/cpuregs/regs[9][2] ;
 wire \soc/cpu/cpuregs/regs[9][30] ;
 wire \soc/cpu/cpuregs/regs[9][31] ;
 wire \soc/cpu/cpuregs/regs[9][3] ;
 wire \soc/cpu/cpuregs/regs[9][4] ;
 wire \soc/cpu/cpuregs/regs[9][5] ;
 wire \soc/cpu/cpuregs/regs[9][6] ;
 wire \soc/cpu/cpuregs/regs[9][7] ;
 wire \soc/cpu/cpuregs/regs[9][8] ;
 wire \soc/cpu/cpuregs/regs[9][9] ;
 wire \soc/simpleuart/_0000_ ;
 wire \soc/simpleuart/_0001_ ;
 wire \soc/simpleuart/_0002_ ;
 wire \soc/simpleuart/_0003_ ;
 wire \soc/simpleuart/_0004_ ;
 wire \soc/simpleuart/_0005_ ;
 wire \soc/simpleuart/_0006_ ;
 wire \soc/simpleuart/_0007_ ;
 wire \soc/simpleuart/_0008_ ;
 wire \soc/simpleuart/_0009_ ;
 wire \soc/simpleuart/_0010_ ;
 wire \soc/simpleuart/_0011_ ;
 wire \soc/simpleuart/_0012_ ;
 wire \soc/simpleuart/_0013_ ;
 wire \soc/simpleuart/_0014_ ;
 wire \soc/simpleuart/_0015_ ;
 wire \soc/simpleuart/_0016_ ;
 wire \soc/simpleuart/_0017_ ;
 wire \soc/simpleuart/_0018_ ;
 wire \soc/simpleuart/_0019_ ;
 wire \soc/simpleuart/_0020_ ;
 wire \soc/simpleuart/_0021_ ;
 wire \soc/simpleuart/_0022_ ;
 wire \soc/simpleuart/_0023_ ;
 wire \soc/simpleuart/_0024_ ;
 wire \soc/simpleuart/_0025_ ;
 wire \soc/simpleuart/_0026_ ;
 wire \soc/simpleuart/_0027_ ;
 wire \soc/simpleuart/_0028_ ;
 wire \soc/simpleuart/_0029_ ;
 wire \soc/simpleuart/_0030_ ;
 wire \soc/simpleuart/_0031_ ;
 wire \soc/simpleuart/_0032_ ;
 wire \soc/simpleuart/_0033_ ;
 wire \soc/simpleuart/_0034_ ;
 wire \soc/simpleuart/_0035_ ;
 wire \soc/simpleuart/_0036_ ;
 wire \soc/simpleuart/_0037_ ;
 wire \soc/simpleuart/_0038_ ;
 wire \soc/simpleuart/_0039_ ;
 wire \soc/simpleuart/_0040_ ;
 wire \soc/simpleuart/_0041_ ;
 wire \soc/simpleuart/_0042_ ;
 wire \soc/simpleuart/_0043_ ;
 wire \soc/simpleuart/_0044_ ;
 wire \soc/simpleuart/_0045_ ;
 wire \soc/simpleuart/_0046_ ;
 wire \soc/simpleuart/_0047_ ;
 wire \soc/simpleuart/_0048_ ;
 wire \soc/simpleuart/_0049_ ;
 wire \soc/simpleuart/_0050_ ;
 wire \soc/simpleuart/_0051_ ;
 wire \soc/simpleuart/_0052_ ;
 wire \soc/simpleuart/_0053_ ;
 wire \soc/simpleuart/_0054_ ;
 wire \soc/simpleuart/_0055_ ;
 wire \soc/simpleuart/_0056_ ;
 wire \soc/simpleuart/_0057_ ;
 wire \soc/simpleuart/_0058_ ;
 wire \soc/simpleuart/_0059_ ;
 wire \soc/simpleuart/_0060_ ;
 wire \soc/simpleuart/_0061_ ;
 wire \soc/simpleuart/_0062_ ;
 wire \soc/simpleuart/_0063_ ;
 wire \soc/simpleuart/_0064_ ;
 wire \soc/simpleuart/_0065_ ;
 wire \soc/simpleuart/_0066_ ;
 wire \soc/simpleuart/_0067_ ;
 wire \soc/simpleuart/_0068_ ;
 wire \soc/simpleuart/_0069_ ;
 wire \soc/simpleuart/_0070_ ;
 wire \soc/simpleuart/_0071_ ;
 wire \soc/simpleuart/_0072_ ;
 wire \soc/simpleuart/_0073_ ;
 wire \soc/simpleuart/_0074_ ;
 wire \soc/simpleuart/_0075_ ;
 wire \soc/simpleuart/_0076_ ;
 wire \soc/simpleuart/_0077_ ;
 wire \soc/simpleuart/_0078_ ;
 wire \soc/simpleuart/_0079_ ;
 wire \soc/simpleuart/_0080_ ;
 wire \soc/simpleuart/_0081_ ;
 wire \soc/simpleuart/_0082_ ;
 wire \soc/simpleuart/_0083_ ;
 wire \soc/simpleuart/_0084_ ;
 wire \soc/simpleuart/_0085_ ;
 wire \soc/simpleuart/_0086_ ;
 wire \soc/simpleuart/_0087_ ;
 wire \soc/simpleuart/_0088_ ;
 wire \soc/simpleuart/_0089_ ;
 wire \soc/simpleuart/_0090_ ;
 wire \soc/simpleuart/_0091_ ;
 wire \soc/simpleuart/_0092_ ;
 wire \soc/simpleuart/_0093_ ;
 wire \soc/simpleuart/_0094_ ;
 wire \soc/simpleuart/_0095_ ;
 wire \soc/simpleuart/_0096_ ;
 wire \soc/simpleuart/_0097_ ;
 wire \soc/simpleuart/_0098_ ;
 wire \soc/simpleuart/_0099_ ;
 wire \soc/simpleuart/_0100_ ;
 wire \soc/simpleuart/_0101_ ;
 wire \soc/simpleuart/_0102_ ;
 wire \soc/simpleuart/_0103_ ;
 wire \soc/simpleuart/_0104_ ;
 wire \soc/simpleuart/_0105_ ;
 wire \soc/simpleuart/_0106_ ;
 wire \soc/simpleuart/_0107_ ;
 wire \soc/simpleuart/_0108_ ;
 wire \soc/simpleuart/_0109_ ;
 wire \soc/simpleuart/_0110_ ;
 wire \soc/simpleuart/_0111_ ;
 wire \soc/simpleuart/_0112_ ;
 wire \soc/simpleuart/_0113_ ;
 wire \soc/simpleuart/_0114_ ;
 wire \soc/simpleuart/_0115_ ;
 wire \soc/simpleuart/_0116_ ;
 wire \soc/simpleuart/_0117_ ;
 wire \soc/simpleuart/_0118_ ;
 wire \soc/simpleuart/_0119_ ;
 wire \soc/simpleuart/_0120_ ;
 wire \soc/simpleuart/_0121_ ;
 wire \soc/simpleuart/_0122_ ;
 wire \soc/simpleuart/_0123_ ;
 wire \soc/simpleuart/_0124_ ;
 wire \soc/simpleuart/_0125_ ;
 wire \soc/simpleuart/_0126_ ;
 wire \soc/simpleuart/_0127_ ;
 wire \soc/simpleuart/_0128_ ;
 wire \soc/simpleuart/_0129_ ;
 wire \soc/simpleuart/_0130_ ;
 wire \soc/simpleuart/_0131_ ;
 wire \soc/simpleuart/_0132_ ;
 wire \soc/simpleuart/_0133_ ;
 wire \soc/simpleuart/_0134_ ;
 wire net346;
 wire \soc/simpleuart/_0136_ ;
 wire \soc/simpleuart/_0137_ ;
 wire \soc/simpleuart/_0138_ ;
 wire \soc/simpleuart/_0139_ ;
 wire \soc/simpleuart/_0140_ ;
 wire \soc/simpleuart/_0141_ ;
 wire \soc/simpleuart/_0142_ ;
 wire \soc/simpleuart/_0143_ ;
 wire \soc/simpleuart/_0144_ ;
 wire \soc/simpleuart/_0145_ ;
 wire \soc/simpleuart/_0146_ ;
 wire \soc/simpleuart/_0147_ ;
 wire \soc/simpleuart/_0148_ ;
 wire \soc/simpleuart/_0149_ ;
 wire \soc/simpleuart/_0150_ ;
 wire \soc/simpleuart/_0151_ ;
 wire \soc/simpleuart/_0152_ ;
 wire \soc/simpleuart/_0153_ ;
 wire \soc/simpleuart/_0154_ ;
 wire \soc/simpleuart/_0155_ ;
 wire \soc/simpleuart/_0156_ ;
 wire \soc/simpleuart/_0157_ ;
 wire \soc/simpleuart/_0158_ ;
 wire \soc/simpleuart/_0159_ ;
 wire \soc/simpleuart/_0160_ ;
 wire \soc/simpleuart/_0161_ ;
 wire \soc/simpleuart/_0162_ ;
 wire \soc/simpleuart/_0163_ ;
 wire \soc/simpleuart/_0164_ ;
 wire \soc/simpleuart/_0165_ ;
 wire \soc/simpleuart/_0166_ ;
 wire \soc/simpleuart/_0167_ ;
 wire \soc/simpleuart/_0168_ ;
 wire \soc/simpleuart/_0169_ ;
 wire \soc/simpleuart/_0170_ ;
 wire \soc/simpleuart/_0171_ ;
 wire \soc/simpleuart/_0172_ ;
 wire \soc/simpleuart/_0173_ ;
 wire \soc/simpleuart/_0174_ ;
 wire \soc/simpleuart/_0175_ ;
 wire \soc/simpleuart/_0176_ ;
 wire \soc/simpleuart/_0177_ ;
 wire \soc/simpleuart/_0178_ ;
 wire \soc/simpleuart/_0179_ ;
 wire \soc/simpleuart/_0180_ ;
 wire \soc/simpleuart/_0181_ ;
 wire \soc/simpleuart/_0182_ ;
 wire \soc/simpleuart/_0183_ ;
 wire \soc/simpleuart/_0184_ ;
 wire \soc/simpleuart/_0185_ ;
 wire \soc/simpleuart/_0186_ ;
 wire \soc/simpleuart/_0187_ ;
 wire \soc/simpleuart/_0188_ ;
 wire \soc/simpleuart/_0189_ ;
 wire \soc/simpleuart/_0190_ ;
 wire \soc/simpleuart/_0191_ ;
 wire \soc/simpleuart/_0192_ ;
 wire \soc/simpleuart/_0193_ ;
 wire \soc/simpleuart/_0194_ ;
 wire \soc/simpleuart/_0195_ ;
 wire \soc/simpleuart/_0196_ ;
 wire \soc/simpleuart/_0197_ ;
 wire \soc/simpleuart/_0198_ ;
 wire \soc/simpleuart/_0199_ ;
 wire \soc/simpleuart/_0200_ ;
 wire \soc/simpleuart/_0201_ ;
 wire \soc/simpleuart/_0202_ ;
 wire \soc/simpleuart/_0203_ ;
 wire \soc/simpleuart/_0204_ ;
 wire \soc/simpleuart/_0205_ ;
 wire \soc/simpleuart/_0206_ ;
 wire \soc/simpleuart/_0207_ ;
 wire \soc/simpleuart/_0208_ ;
 wire \soc/simpleuart/_0209_ ;
 wire \soc/simpleuart/_0210_ ;
 wire \soc/simpleuart/_0211_ ;
 wire \soc/simpleuart/_0212_ ;
 wire \soc/simpleuart/_0213_ ;
 wire \soc/simpleuart/_0214_ ;
 wire \soc/simpleuart/_0215_ ;
 wire \soc/simpleuart/_0216_ ;
 wire \soc/simpleuart/_0217_ ;
 wire \soc/simpleuart/_0218_ ;
 wire \soc/simpleuart/_0219_ ;
 wire \soc/simpleuart/_0220_ ;
 wire \soc/simpleuart/_0221_ ;
 wire \soc/simpleuart/_0222_ ;
 wire net345;
 wire \soc/simpleuart/_0224_ ;
 wire \soc/simpleuart/_0225_ ;
 wire \soc/simpleuart/_0226_ ;
 wire \soc/simpleuart/_0227_ ;
 wire \soc/simpleuart/_0228_ ;
 wire \soc/simpleuart/_0229_ ;
 wire \soc/simpleuart/_0230_ ;
 wire \soc/simpleuart/_0231_ ;
 wire \soc/simpleuart/_0232_ ;
 wire \soc/simpleuart/_0233_ ;
 wire \soc/simpleuart/_0234_ ;
 wire \soc/simpleuart/_0235_ ;
 wire \soc/simpleuart/_0236_ ;
 wire \soc/simpleuart/_0237_ ;
 wire \soc/simpleuart/_0238_ ;
 wire \soc/simpleuart/_0239_ ;
 wire \soc/simpleuart/_0240_ ;
 wire \soc/simpleuart/_0241_ ;
 wire \soc/simpleuart/_0242_ ;
 wire \soc/simpleuart/_0243_ ;
 wire \soc/simpleuart/_0244_ ;
 wire \soc/simpleuart/_0245_ ;
 wire \soc/simpleuart/_0246_ ;
 wire \soc/simpleuart/_0247_ ;
 wire \soc/simpleuart/_0248_ ;
 wire \soc/simpleuart/_0249_ ;
 wire \soc/simpleuart/_0250_ ;
 wire \soc/simpleuart/_0251_ ;
 wire \soc/simpleuart/_0252_ ;
 wire \soc/simpleuart/_0253_ ;
 wire \soc/simpleuart/_0254_ ;
 wire \soc/simpleuart/_0255_ ;
 wire \soc/simpleuart/_0256_ ;
 wire net344;
 wire \soc/simpleuart/_0258_ ;
 wire \soc/simpleuart/_0259_ ;
 wire net343;
 wire \soc/simpleuart/_0261_ ;
 wire \soc/simpleuart/_0262_ ;
 wire \soc/simpleuart/_0263_ ;
 wire net342;
 wire \soc/simpleuart/_0265_ ;
 wire \soc/simpleuart/_0266_ ;
 wire \soc/simpleuart/_0267_ ;
 wire \soc/simpleuart/_0268_ ;
 wire \soc/simpleuart/_0269_ ;
 wire \soc/simpleuart/_0270_ ;
 wire \soc/simpleuart/_0271_ ;
 wire \soc/simpleuart/_0272_ ;
 wire \soc/simpleuart/_0273_ ;
 wire \soc/simpleuart/_0274_ ;
 wire \soc/simpleuart/_0275_ ;
 wire \soc/simpleuart/_0276_ ;
 wire \soc/simpleuart/_0277_ ;
 wire \soc/simpleuart/_0278_ ;
 wire \soc/simpleuart/_0279_ ;
 wire \soc/simpleuart/_0280_ ;
 wire net341;
 wire \soc/simpleuart/_0282_ ;
 wire net340;
 wire \soc/simpleuart/_0284_ ;
 wire \soc/simpleuart/_0285_ ;
 wire \soc/simpleuart/_0286_ ;
 wire \soc/simpleuart/_0287_ ;
 wire \soc/simpleuart/_0288_ ;
 wire \soc/simpleuart/_0289_ ;
 wire \soc/simpleuart/_0290_ ;
 wire \soc/simpleuart/_0291_ ;
 wire \soc/simpleuart/_0292_ ;
 wire \soc/simpleuart/_0293_ ;
 wire \soc/simpleuart/_0294_ ;
 wire \soc/simpleuart/_0295_ ;
 wire \soc/simpleuart/_0296_ ;
 wire \soc/simpleuart/_0297_ ;
 wire \soc/simpleuart/_0298_ ;
 wire \soc/simpleuart/_0299_ ;
 wire \soc/simpleuart/_0300_ ;
 wire \soc/simpleuart/_0301_ ;
 wire \soc/simpleuart/_0302_ ;
 wire \soc/simpleuart/_0303_ ;
 wire \soc/simpleuart/_0304_ ;
 wire \soc/simpleuart/_0305_ ;
 wire net339;
 wire \soc/simpleuart/_0307_ ;
 wire \soc/simpleuart/_0308_ ;
 wire \soc/simpleuart/_0309_ ;
 wire \soc/simpleuart/_0310_ ;
 wire \soc/simpleuart/_0311_ ;
 wire \soc/simpleuart/_0312_ ;
 wire \soc/simpleuart/_0313_ ;
 wire \soc/simpleuart/_0314_ ;
 wire \soc/simpleuart/_0315_ ;
 wire \soc/simpleuart/_0316_ ;
 wire \soc/simpleuart/_0317_ ;
 wire \soc/simpleuart/_0318_ ;
 wire \soc/simpleuart/_0319_ ;
 wire \soc/simpleuart/_0320_ ;
 wire \soc/simpleuart/_0321_ ;
 wire \soc/simpleuart/_0322_ ;
 wire \soc/simpleuart/_0323_ ;
 wire \soc/simpleuart/_0324_ ;
 wire \soc/simpleuart/_0325_ ;
 wire \soc/simpleuart/_0326_ ;
 wire \soc/simpleuart/_0327_ ;
 wire \soc/simpleuart/_0328_ ;
 wire \soc/simpleuart/_0329_ ;
 wire \soc/simpleuart/_0330_ ;
 wire \soc/simpleuart/_0331_ ;
 wire \soc/simpleuart/_0332_ ;
 wire \soc/simpleuart/_0333_ ;
 wire \soc/simpleuart/_0334_ ;
 wire \soc/simpleuart/_0335_ ;
 wire \soc/simpleuart/_0336_ ;
 wire net338;
 wire \soc/simpleuart/_0338_ ;
 wire \soc/simpleuart/_0339_ ;
 wire net337;
 wire net336;
 wire \soc/simpleuart/_0342_ ;
 wire \soc/simpleuart/_0343_ ;
 wire \soc/simpleuart/_0344_ ;
 wire \soc/simpleuart/_0345_ ;
 wire \soc/simpleuart/_0346_ ;
 wire \soc/simpleuart/_0347_ ;
 wire \soc/simpleuart/_0348_ ;
 wire \soc/simpleuart/_0349_ ;
 wire \soc/simpleuart/_0350_ ;
 wire \soc/simpleuart/_0351_ ;
 wire \soc/simpleuart/_0352_ ;
 wire \soc/simpleuart/_0353_ ;
 wire net335;
 wire \soc/simpleuart/_0355_ ;
 wire \soc/simpleuart/_0356_ ;
 wire \soc/simpleuart/_0357_ ;
 wire \soc/simpleuart/_0358_ ;
 wire \soc/simpleuart/_0359_ ;
 wire \soc/simpleuart/_0360_ ;
 wire net334;
 wire \soc/simpleuart/_0362_ ;
 wire \soc/simpleuart/_0363_ ;
 wire \soc/simpleuart/_0364_ ;
 wire \soc/simpleuart/_0365_ ;
 wire \soc/simpleuart/_0366_ ;
 wire \soc/simpleuart/_0367_ ;
 wire net333;
 wire \soc/simpleuart/_0369_ ;
 wire \soc/simpleuart/_0370_ ;
 wire \soc/simpleuart/_0371_ ;
 wire \soc/simpleuart/_0372_ ;
 wire \soc/simpleuart/_0373_ ;
 wire \soc/simpleuart/_0374_ ;
 wire \soc/simpleuart/_0375_ ;
 wire \soc/simpleuart/_0376_ ;
 wire \soc/simpleuart/_0377_ ;
 wire net332;
 wire \soc/simpleuart/_0379_ ;
 wire \soc/simpleuart/_0380_ ;
 wire \soc/simpleuart/_0381_ ;
 wire \soc/simpleuart/_0382_ ;
 wire \soc/simpleuart/_0383_ ;
 wire \soc/simpleuart/_0384_ ;
 wire \soc/simpleuart/_0385_ ;
 wire \soc/simpleuart/_0386_ ;
 wire \soc/simpleuart/_0387_ ;
 wire \soc/simpleuart/_0388_ ;
 wire \soc/simpleuart/_0389_ ;
 wire \soc/simpleuart/_0390_ ;
 wire \soc/simpleuart/_0391_ ;
 wire \soc/simpleuart/_0392_ ;
 wire \soc/simpleuart/_0393_ ;
 wire \soc/simpleuart/_0394_ ;
 wire \soc/simpleuart/_0395_ ;
 wire \soc/simpleuart/_0396_ ;
 wire \soc/simpleuart/_0397_ ;
 wire \soc/simpleuart/_0398_ ;
 wire \soc/simpleuart/_0399_ ;
 wire \soc/simpleuart/_0400_ ;
 wire \soc/simpleuart/_0401_ ;
 wire \soc/simpleuart/_0402_ ;
 wire \soc/simpleuart/_0403_ ;
 wire \soc/simpleuart/_0404_ ;
 wire \soc/simpleuart/_0405_ ;
 wire \soc/simpleuart/_0406_ ;
 wire \soc/simpleuart/_0407_ ;
 wire \soc/simpleuart/_0408_ ;
 wire \soc/simpleuart/_0409_ ;
 wire \soc/simpleuart/_0410_ ;
 wire \soc/simpleuart/_0411_ ;
 wire \soc/simpleuart/_0412_ ;
 wire net331;
 wire \soc/simpleuart/_0414_ ;
 wire \soc/simpleuart/_0415_ ;
 wire \soc/simpleuart/_0416_ ;
 wire net330;
 wire \soc/simpleuart/_0418_ ;
 wire \soc/simpleuart/_0419_ ;
 wire \soc/simpleuart/_0420_ ;
 wire \soc/simpleuart/_0421_ ;
 wire \soc/simpleuart/_0422_ ;
 wire \soc/simpleuart/_0423_ ;
 wire \soc/simpleuart/_0424_ ;
 wire \soc/simpleuart/_0425_ ;
 wire \soc/simpleuart/_0426_ ;
 wire \soc/simpleuart/_0427_ ;
 wire \soc/simpleuart/_0428_ ;
 wire \soc/simpleuart/_0429_ ;
 wire \soc/simpleuart/_0430_ ;
 wire \soc/simpleuart/_0431_ ;
 wire \soc/simpleuart/_0432_ ;
 wire \soc/simpleuart/_0433_ ;
 wire \soc/simpleuart/_0434_ ;
 wire \soc/simpleuart/_0435_ ;
 wire \soc/simpleuart/_0436_ ;
 wire \soc/simpleuart/_0437_ ;
 wire \soc/simpleuart/_0438_ ;
 wire \soc/simpleuart/_0439_ ;
 wire \soc/simpleuart/_0440_ ;
 wire \soc/simpleuart/_0441_ ;
 wire \soc/simpleuart/_0442_ ;
 wire \soc/simpleuart/_0443_ ;
 wire \soc/simpleuart/_0444_ ;
 wire \soc/simpleuart/_0445_ ;
 wire \soc/simpleuart/_0446_ ;
 wire \soc/simpleuart/_0447_ ;
 wire \soc/simpleuart/_0448_ ;
 wire \soc/simpleuart/_0449_ ;
 wire \soc/simpleuart/_0450_ ;
 wire \soc/simpleuart/_0451_ ;
 wire \soc/simpleuart/_0452_ ;
 wire \soc/simpleuart/_0453_ ;
 wire \soc/simpleuart/_0454_ ;
 wire \soc/simpleuart/_0455_ ;
 wire \soc/simpleuart/_0456_ ;
 wire \soc/simpleuart/_0457_ ;
 wire \soc/simpleuart/_0458_ ;
 wire \soc/simpleuart/_0459_ ;
 wire \soc/simpleuart/_0460_ ;
 wire \soc/simpleuart/_0461_ ;
 wire \soc/simpleuart/_0462_ ;
 wire \soc/simpleuart/_0463_ ;
 wire \soc/simpleuart/_0464_ ;
 wire \soc/simpleuart/_0465_ ;
 wire \soc/simpleuart/_0466_ ;
 wire \soc/simpleuart/_0467_ ;
 wire \soc/simpleuart/_0468_ ;
 wire \soc/simpleuart/_0469_ ;
 wire \soc/simpleuart/_0470_ ;
 wire \soc/simpleuart/_0471_ ;
 wire \soc/simpleuart/_0472_ ;
 wire \soc/simpleuart/_0473_ ;
 wire \soc/simpleuart/_0474_ ;
 wire \soc/simpleuart/_0475_ ;
 wire \soc/simpleuart/_0476_ ;
 wire \soc/simpleuart/_0477_ ;
 wire \soc/simpleuart/_0478_ ;
 wire \soc/simpleuart/_0479_ ;
 wire \soc/simpleuart/_0480_ ;
 wire \soc/simpleuart/_0481_ ;
 wire \soc/simpleuart/_0482_ ;
 wire \soc/simpleuart/_0483_ ;
 wire \soc/simpleuart/_0484_ ;
 wire \soc/simpleuart/_0485_ ;
 wire \soc/simpleuart/_0486_ ;
 wire \soc/simpleuart/_0487_ ;
 wire \soc/simpleuart/_0488_ ;
 wire \soc/simpleuart/_0489_ ;
 wire \soc/simpleuart/_0490_ ;
 wire \soc/simpleuart/_0491_ ;
 wire \soc/simpleuart/_0492_ ;
 wire \soc/simpleuart/_0493_ ;
 wire \soc/simpleuart/_0494_ ;
 wire \soc/simpleuart/_0495_ ;
 wire \soc/simpleuart/_0496_ ;
 wire \soc/simpleuart/_0497_ ;
 wire \soc/simpleuart/_0498_ ;
 wire \soc/simpleuart/_0499_ ;
 wire \soc/simpleuart/_0500_ ;
 wire \soc/simpleuart/_0501_ ;
 wire \soc/simpleuart/_0502_ ;
 wire \soc/simpleuart/_0503_ ;
 wire \soc/simpleuart/_0504_ ;
 wire \soc/simpleuart/_0505_ ;
 wire \soc/simpleuart/_0506_ ;
 wire \soc/simpleuart/_0507_ ;
 wire \soc/simpleuart/_0508_ ;
 wire \soc/simpleuart/_0509_ ;
 wire \soc/simpleuart/_0510_ ;
 wire \soc/simpleuart/_0511_ ;
 wire \soc/simpleuart/_0512_ ;
 wire \soc/simpleuart/_0513_ ;
 wire \soc/simpleuart/_0514_ ;
 wire \soc/simpleuart/_0515_ ;
 wire \soc/simpleuart/_0516_ ;
 wire \soc/simpleuart/_0517_ ;
 wire \soc/simpleuart/_0518_ ;
 wire \soc/simpleuart/_0519_ ;
 wire \soc/simpleuart/_0520_ ;
 wire \soc/simpleuart/_0521_ ;
 wire \soc/simpleuart/_0522_ ;
 wire \soc/simpleuart/_0523_ ;
 wire \soc/simpleuart/_0524_ ;
 wire \soc/simpleuart/_0525_ ;
 wire \soc/simpleuart/_0526_ ;
 wire \soc/simpleuart/_0527_ ;
 wire \soc/simpleuart/_0528_ ;
 wire \soc/simpleuart/_0529_ ;
 wire \soc/simpleuart/_0530_ ;
 wire \soc/simpleuart/_0531_ ;
 wire \soc/simpleuart/_0532_ ;
 wire \soc/simpleuart/_0533_ ;
 wire \soc/simpleuart/_0534_ ;
 wire \soc/simpleuart/_0535_ ;
 wire \soc/simpleuart/_0536_ ;
 wire \soc/simpleuart/_0537_ ;
 wire \soc/simpleuart/_0538_ ;
 wire \soc/simpleuart/_0539_ ;
 wire \soc/simpleuart/_0540_ ;
 wire \soc/simpleuart/_0541_ ;
 wire \soc/simpleuart/_0542_ ;
 wire \soc/simpleuart/_0543_ ;
 wire \soc/simpleuart/_0544_ ;
 wire \soc/simpleuart/_0545_ ;
 wire \soc/simpleuart/_0546_ ;
 wire \soc/simpleuart/_0547_ ;
 wire \soc/simpleuart/_0548_ ;
 wire \soc/simpleuart/_0549_ ;
 wire \soc/simpleuart/_0550_ ;
 wire \soc/simpleuart/_0551_ ;
 wire \soc/simpleuart/_0552_ ;
 wire \soc/simpleuart/_0553_ ;
 wire \soc/simpleuart/_0554_ ;
 wire \soc/simpleuart/_0555_ ;
 wire \soc/simpleuart/_0556_ ;
 wire \soc/simpleuart/_0557_ ;
 wire \soc/simpleuart/_0558_ ;
 wire \soc/simpleuart/_0559_ ;
 wire \soc/simpleuart/_0560_ ;
 wire \soc/simpleuart/_0561_ ;
 wire \soc/simpleuart/_0562_ ;
 wire \soc/simpleuart/_0563_ ;
 wire \soc/simpleuart/_0564_ ;
 wire \soc/simpleuart/_0565_ ;
 wire \soc/simpleuart/_0566_ ;
 wire \soc/simpleuart/_0567_ ;
 wire \soc/simpleuart/_0568_ ;
 wire \soc/simpleuart/_0569_ ;
 wire \soc/simpleuart/_0570_ ;
 wire \soc/simpleuart/_0571_ ;
 wire \soc/simpleuart/_0572_ ;
 wire \soc/simpleuart/_0573_ ;
 wire \soc/simpleuart/_0574_ ;
 wire \soc/simpleuart/_0575_ ;
 wire \soc/simpleuart/_0576_ ;
 wire \soc/simpleuart/_0577_ ;
 wire \soc/simpleuart/_0578_ ;
 wire \soc/simpleuart/_0579_ ;
 wire net329;
 wire \soc/simpleuart/_0581_ ;
 wire \soc/simpleuart/_0582_ ;
 wire \soc/simpleuart/_0583_ ;
 wire \soc/simpleuart/_0584_ ;
 wire \soc/simpleuart/_0585_ ;
 wire \soc/simpleuart/_0586_ ;
 wire \soc/simpleuart/_0587_ ;
 wire \soc/simpleuart/_0588_ ;
 wire \soc/simpleuart/_0589_ ;
 wire \soc/simpleuart/_0590_ ;
 wire \soc/simpleuart/_0591_ ;
 wire \soc/simpleuart/_0592_ ;
 wire \soc/simpleuart/_0593_ ;
 wire \soc/simpleuart/_0594_ ;
 wire \soc/simpleuart/_0595_ ;
 wire \soc/simpleuart/_0596_ ;
 wire net328;
 wire net327;
 wire \soc/simpleuart/_0599_ ;
 wire \soc/simpleuart/_0600_ ;
 wire \soc/simpleuart/_0601_ ;
 wire \soc/simpleuart/_0602_ ;
 wire \soc/simpleuart/_0603_ ;
 wire \soc/simpleuart/_0604_ ;
 wire \soc/simpleuart/_0605_ ;
 wire \soc/simpleuart/_0606_ ;
 wire \soc/simpleuart/_0607_ ;
 wire net326;
 wire \soc/simpleuart/_0609_ ;
 wire net325;
 wire \soc/simpleuart/_0611_ ;
 wire \soc/simpleuart/_0612_ ;
 wire \soc/simpleuart/_0613_ ;
 wire \soc/simpleuart/_0614_ ;
 wire \soc/simpleuart/_0615_ ;
 wire \soc/simpleuart/_0616_ ;
 wire \soc/simpleuart/_0617_ ;
 wire net324;
 wire \soc/simpleuart/_0619_ ;
 wire \soc/simpleuart/_0620_ ;
 wire \soc/simpleuart/_0621_ ;
 wire \soc/simpleuart/_0622_ ;
 wire \soc/simpleuart/_0623_ ;
 wire \soc/simpleuart/_0624_ ;
 wire \soc/simpleuart/_0625_ ;
 wire \soc/simpleuart/_0626_ ;
 wire \soc/simpleuart/_0627_ ;
 wire \soc/simpleuart/_0628_ ;
 wire \soc/simpleuart/_0629_ ;
 wire \soc/simpleuart/_0630_ ;
 wire \soc/simpleuart/_0631_ ;
 wire \soc/simpleuart/_0632_ ;
 wire \soc/simpleuart/_0633_ ;
 wire \soc/simpleuart/_0634_ ;
 wire \soc/simpleuart/_0635_ ;
 wire \soc/simpleuart/_0636_ ;
 wire \soc/simpleuart/_0637_ ;
 wire \soc/simpleuart/_0638_ ;
 wire \soc/simpleuart/_0639_ ;
 wire \soc/simpleuart/_0640_ ;
 wire \soc/simpleuart/_0641_ ;
 wire \soc/simpleuart/_0642_ ;
 wire \soc/simpleuart/_0643_ ;
 wire \soc/simpleuart/_0644_ ;
 wire \soc/simpleuart/_0645_ ;
 wire \soc/simpleuart/_0646_ ;
 wire \soc/simpleuart/_0647_ ;
 wire \soc/simpleuart/_0648_ ;
 wire \soc/simpleuart/_0649_ ;
 wire \soc/simpleuart/_0650_ ;
 wire \soc/simpleuart/_0651_ ;
 wire \soc/simpleuart/_0652_ ;
 wire \soc/simpleuart/_0653_ ;
 wire \soc/simpleuart/_0654_ ;
 wire \soc/simpleuart/_0655_ ;
 wire \soc/simpleuart/_0656_ ;
 wire \soc/simpleuart/_0657_ ;
 wire \soc/simpleuart/_0658_ ;
 wire \soc/simpleuart/_0659_ ;
 wire \soc/simpleuart/_0660_ ;
 wire \soc/simpleuart/_0661_ ;
 wire \soc/simpleuart/_0662_ ;
 wire \soc/simpleuart/_0663_ ;
 wire net323;
 wire \soc/simpleuart/_0665_ ;
 wire \soc/simpleuart/_0666_ ;
 wire \soc/simpleuart/_0667_ ;
 wire \soc/simpleuart/_0668_ ;
 wire \soc/simpleuart/_0669_ ;
 wire \soc/simpleuart/_0670_ ;
 wire \soc/simpleuart/_0671_ ;
 wire \soc/simpleuart/_0672_ ;
 wire \soc/simpleuart/recv_buf_data[0] ;
 wire \soc/simpleuart/recv_buf_data[1] ;
 wire \soc/simpleuart/recv_buf_data[2] ;
 wire \soc/simpleuart/recv_buf_data[3] ;
 wire \soc/simpleuart/recv_buf_data[4] ;
 wire \soc/simpleuart/recv_buf_data[5] ;
 wire \soc/simpleuart/recv_buf_data[6] ;
 wire \soc/simpleuart/recv_buf_data[7] ;
 wire \soc/simpleuart/recv_buf_valid ;
 wire \soc/simpleuart/recv_divcnt[0] ;
 wire \soc/simpleuart/recv_divcnt[10] ;
 wire \soc/simpleuart/recv_divcnt[11] ;
 wire \soc/simpleuart/recv_divcnt[12] ;
 wire \soc/simpleuart/recv_divcnt[13] ;
 wire \soc/simpleuart/recv_divcnt[14] ;
 wire \soc/simpleuart/recv_divcnt[15] ;
 wire \soc/simpleuart/recv_divcnt[16] ;
 wire \soc/simpleuart/recv_divcnt[17] ;
 wire \soc/simpleuart/recv_divcnt[18] ;
 wire \soc/simpleuart/recv_divcnt[19] ;
 wire \soc/simpleuart/recv_divcnt[1] ;
 wire \soc/simpleuart/recv_divcnt[20] ;
 wire \soc/simpleuart/recv_divcnt[21] ;
 wire \soc/simpleuart/recv_divcnt[22] ;
 wire \soc/simpleuart/recv_divcnt[23] ;
 wire \soc/simpleuart/recv_divcnt[24] ;
 wire \soc/simpleuart/recv_divcnt[25] ;
 wire \soc/simpleuart/recv_divcnt[26] ;
 wire \soc/simpleuart/recv_divcnt[27] ;
 wire \soc/simpleuart/recv_divcnt[28] ;
 wire \soc/simpleuart/recv_divcnt[29] ;
 wire \soc/simpleuart/recv_divcnt[2] ;
 wire \soc/simpleuart/recv_divcnt[30] ;
 wire \soc/simpleuart/recv_divcnt[31] ;
 wire \soc/simpleuart/recv_divcnt[3] ;
 wire \soc/simpleuart/recv_divcnt[4] ;
 wire \soc/simpleuart/recv_divcnt[5] ;
 wire \soc/simpleuart/recv_divcnt[6] ;
 wire \soc/simpleuart/recv_divcnt[7] ;
 wire \soc/simpleuart/recv_divcnt[8] ;
 wire \soc/simpleuart/recv_divcnt[9] ;
 wire \soc/simpleuart/recv_pattern[0] ;
 wire \soc/simpleuart/recv_pattern[1] ;
 wire \soc/simpleuart/recv_pattern[2] ;
 wire \soc/simpleuart/recv_pattern[3] ;
 wire \soc/simpleuart/recv_pattern[4] ;
 wire \soc/simpleuart/recv_pattern[5] ;
 wire \soc/simpleuart/recv_pattern[6] ;
 wire \soc/simpleuart/recv_pattern[7] ;
 wire \soc/simpleuart/recv_state[0] ;
 wire \soc/simpleuart/recv_state[1] ;
 wire \soc/simpleuart/recv_state[2] ;
 wire \soc/simpleuart/recv_state[3] ;
 wire \soc/simpleuart/send_bitcnt[0] ;
 wire \soc/simpleuart/send_bitcnt[1] ;
 wire \soc/simpleuart/send_bitcnt[2] ;
 wire \soc/simpleuart/send_bitcnt[3] ;
 wire \soc/simpleuart/send_divcnt[0] ;
 wire \soc/simpleuart/send_divcnt[10] ;
 wire \soc/simpleuart/send_divcnt[11] ;
 wire \soc/simpleuart/send_divcnt[12] ;
 wire \soc/simpleuart/send_divcnt[13] ;
 wire \soc/simpleuart/send_divcnt[14] ;
 wire \soc/simpleuart/send_divcnt[15] ;
 wire \soc/simpleuart/send_divcnt[16] ;
 wire \soc/simpleuart/send_divcnt[17] ;
 wire \soc/simpleuart/send_divcnt[18] ;
 wire \soc/simpleuart/send_divcnt[19] ;
 wire \soc/simpleuart/send_divcnt[1] ;
 wire \soc/simpleuart/send_divcnt[20] ;
 wire \soc/simpleuart/send_divcnt[21] ;
 wire \soc/simpleuart/send_divcnt[22] ;
 wire \soc/simpleuart/send_divcnt[23] ;
 wire \soc/simpleuart/send_divcnt[24] ;
 wire \soc/simpleuart/send_divcnt[25] ;
 wire \soc/simpleuart/send_divcnt[26] ;
 wire \soc/simpleuart/send_divcnt[27] ;
 wire \soc/simpleuart/send_divcnt[28] ;
 wire \soc/simpleuart/send_divcnt[29] ;
 wire \soc/simpleuart/send_divcnt[2] ;
 wire \soc/simpleuart/send_divcnt[30] ;
 wire \soc/simpleuart/send_divcnt[31] ;
 wire \soc/simpleuart/send_divcnt[3] ;
 wire \soc/simpleuart/send_divcnt[4] ;
 wire \soc/simpleuart/send_divcnt[5] ;
 wire \soc/simpleuart/send_divcnt[6] ;
 wire \soc/simpleuart/send_divcnt[7] ;
 wire \soc/simpleuart/send_divcnt[8] ;
 wire \soc/simpleuart/send_divcnt[9] ;
 wire \soc/simpleuart/send_dummy ;
 wire \soc/simpleuart/send_pattern[1] ;
 wire \soc/simpleuart/send_pattern[2] ;
 wire \soc/simpleuart/send_pattern[3] ;
 wire \soc/simpleuart/send_pattern[4] ;
 wire \soc/simpleuart/send_pattern[5] ;
 wire \soc/simpleuart/send_pattern[6] ;
 wire \soc/simpleuart/send_pattern[7] ;
 wire \soc/simpleuart/send_pattern[8] ;
 wire \soc/spimemio/_0000_ ;
 wire \soc/spimemio/_0001_ ;
 wire \soc/spimemio/_0002_ ;
 wire \soc/spimemio/_0003_ ;
 wire \soc/spimemio/_0004_ ;
 wire \soc/spimemio/_0005_ ;
 wire \soc/spimemio/_0006_ ;
 wire \soc/spimemio/_0007_ ;
 wire \soc/spimemio/_0008_ ;
 wire \soc/spimemio/_0009_ ;
 wire \soc/spimemio/_0010_ ;
 wire \soc/spimemio/_0011_ ;
 wire \soc/spimemio/_0012_ ;
 wire clknet_leaf_0_clk;
 wire \soc/spimemio/_0014_ ;
 wire \soc/spimemio/_0015_ ;
 wire \soc/spimemio/_0016_ ;
 wire \soc/spimemio/_0017_ ;
 wire \soc/spimemio/_0018_ ;
 wire \soc/spimemio/_0019_ ;
 wire \soc/spimemio/_0020_ ;
 wire \soc/spimemio/_0021_ ;
 wire \soc/spimemio/_0022_ ;
 wire \soc/spimemio/_0023_ ;
 wire \soc/spimemio/_0024_ ;
 wire \soc/spimemio/_0025_ ;
 wire \soc/spimemio/_0026_ ;
 wire \soc/spimemio/_0027_ ;
 wire \soc/spimemio/_0028_ ;
 wire \soc/spimemio/_0029_ ;
 wire \soc/spimemio/_0030_ ;
 wire \soc/spimemio/_0031_ ;
 wire \soc/spimemio/_0032_ ;
 wire \soc/spimemio/_0033_ ;
 wire \soc/spimemio/_0034_ ;
 wire \soc/spimemio/_0035_ ;
 wire \soc/spimemio/_0036_ ;
 wire \soc/spimemio/_0037_ ;
 wire \soc/spimemio/_0038_ ;
 wire \soc/spimemio/_0039_ ;
 wire \soc/spimemio/_0040_ ;
 wire \soc/spimemio/_0041_ ;
 wire \soc/spimemio/_0042_ ;
 wire \soc/spimemio/_0043_ ;
 wire \soc/spimemio/_0044_ ;
 wire \soc/spimemio/_0045_ ;
 wire \soc/spimemio/_0046_ ;
 wire \soc/spimemio/_0047_ ;
 wire \soc/spimemio/_0048_ ;
 wire \soc/spimemio/_0049_ ;
 wire \soc/spimemio/_0050_ ;
 wire \soc/spimemio/_0051_ ;
 wire \soc/spimemio/_0052_ ;
 wire \soc/spimemio/_0053_ ;
 wire \soc/spimemio/_0054_ ;
 wire \soc/spimemio/_0055_ ;
 wire \soc/spimemio/_0056_ ;
 wire \soc/spimemio/_0057_ ;
 wire \soc/spimemio/_0058_ ;
 wire \soc/spimemio/_0059_ ;
 wire \soc/spimemio/_0060_ ;
 wire \soc/spimemio/_0061_ ;
 wire \soc/spimemio/_0062_ ;
 wire \soc/spimemio/_0063_ ;
 wire \soc/spimemio/_0064_ ;
 wire \soc/spimemio/_0065_ ;
 wire \soc/spimemio/_0066_ ;
 wire \soc/spimemio/_0067_ ;
 wire \soc/spimemio/_0068_ ;
 wire \soc/spimemio/_0069_ ;
 wire \soc/spimemio/_0070_ ;
 wire \soc/spimemio/_0071_ ;
 wire \soc/spimemio/_0072_ ;
 wire \soc/spimemio/_0073_ ;
 wire \soc/spimemio/_0074_ ;
 wire \soc/spimemio/_0075_ ;
 wire \soc/spimemio/_0076_ ;
 wire \soc/spimemio/_0077_ ;
 wire \soc/spimemio/_0078_ ;
 wire \soc/spimemio/_0079_ ;
 wire \soc/spimemio/_0080_ ;
 wire \soc/spimemio/_0081_ ;
 wire \soc/spimemio/_0082_ ;
 wire \soc/spimemio/_0083_ ;
 wire \soc/spimemio/_0084_ ;
 wire \soc/spimemio/_0085_ ;
 wire \soc/spimemio/_0086_ ;
 wire \soc/spimemio/_0087_ ;
 wire \soc/spimemio/_0088_ ;
 wire \soc/spimemio/_0089_ ;
 wire \soc/spimemio/_0090_ ;
 wire \soc/spimemio/_0091_ ;
 wire \soc/spimemio/_0092_ ;
 wire \soc/spimemio/_0093_ ;
 wire \soc/spimemio/_0094_ ;
 wire \soc/spimemio/_0095_ ;
 wire \soc/spimemio/_0096_ ;
 wire \soc/spimemio/_0097_ ;
 wire \soc/spimemio/_0098_ ;
 wire \soc/spimemio/_0099_ ;
 wire \soc/spimemio/_0100_ ;
 wire \soc/spimemio/_0101_ ;
 wire \soc/spimemio/_0102_ ;
 wire \soc/spimemio/_0103_ ;
 wire \soc/spimemio/_0104_ ;
 wire \soc/spimemio/_0105_ ;
 wire \soc/spimemio/_0106_ ;
 wire \soc/spimemio/_0107_ ;
 wire \soc/spimemio/_0108_ ;
 wire \soc/spimemio/_0109_ ;
 wire \soc/spimemio/_0110_ ;
 wire \soc/spimemio/_0111_ ;
 wire \soc/spimemio/_0112_ ;
 wire \soc/spimemio/_0113_ ;
 wire \soc/spimemio/_0114_ ;
 wire \soc/spimemio/_0115_ ;
 wire \soc/spimemio/_0116_ ;
 wire \soc/spimemio/_0117_ ;
 wire \soc/spimemio/_0118_ ;
 wire \soc/spimemio/_0119_ ;
 wire \soc/spimemio/_0120_ ;
 wire \soc/spimemio/_0121_ ;
 wire \soc/spimemio/_0122_ ;
 wire \soc/spimemio/_0123_ ;
 wire \soc/spimemio/_0124_ ;
 wire \soc/spimemio/_0125_ ;
 wire \soc/spimemio/_0126_ ;
 wire \soc/spimemio/_0127_ ;
 wire \soc/spimemio/_0128_ ;
 wire \soc/spimemio/_0129_ ;
 wire \soc/spimemio/_0130_ ;
 wire \soc/spimemio/_0131_ ;
 wire \soc/spimemio/_0132_ ;
 wire \soc/spimemio/_0133_ ;
 wire \soc/spimemio/_0134_ ;
 wire \soc/spimemio/_0135_ ;
 wire \soc/spimemio/_0136_ ;
 wire \soc/spimemio/_0137_ ;
 wire \soc/spimemio/_0138_ ;
 wire \soc/spimemio/_0139_ ;
 wire \soc/spimemio/_0140_ ;
 wire \soc/spimemio/_0141_ ;
 wire net299;
 wire \soc/spimemio/_0143_ ;
 wire \soc/spimemio/_0144_ ;
 wire \soc/spimemio/_0145_ ;
 wire \soc/spimemio/_0146_ ;
 wire \soc/spimemio/_0147_ ;
 wire \soc/spimemio/_0148_ ;
 wire \soc/spimemio/_0149_ ;
 wire \soc/spimemio/_0150_ ;
 wire net298;
 wire \soc/spimemio/_0152_ ;
 wire \soc/spimemio/_0153_ ;
 wire \soc/spimemio/_0154_ ;
 wire \soc/spimemio/_0155_ ;
 wire \soc/spimemio/_0156_ ;
 wire \soc/spimemio/_0157_ ;
 wire \soc/spimemio/_0158_ ;
 wire \soc/spimemio/_0159_ ;
 wire \soc/spimemio/_0160_ ;
 wire \soc/spimemio/_0161_ ;
 wire \soc/spimemio/_0162_ ;
 wire \soc/spimemio/_0163_ ;
 wire \soc/spimemio/_0164_ ;
 wire \soc/spimemio/_0165_ ;
 wire \soc/spimemio/_0166_ ;
 wire \soc/spimemio/_0167_ ;
 wire \soc/spimemio/_0168_ ;
 wire \soc/spimemio/_0169_ ;
 wire \soc/spimemio/_0170_ ;
 wire \soc/spimemio/_0171_ ;
 wire \soc/spimemio/_0172_ ;
 wire \soc/spimemio/_0173_ ;
 wire \soc/spimemio/_0174_ ;
 wire \soc/spimemio/_0175_ ;
 wire \soc/spimemio/_0176_ ;
 wire \soc/spimemio/_0177_ ;
 wire \soc/spimemio/_0178_ ;
 wire \soc/spimemio/_0179_ ;
 wire \soc/spimemio/_0180_ ;
 wire \soc/spimemio/_0181_ ;
 wire \soc/spimemio/_0182_ ;
 wire \soc/spimemio/_0183_ ;
 wire \soc/spimemio/_0184_ ;
 wire net297;
 wire \soc/spimemio/_0186_ ;
 wire net296;
 wire \soc/spimemio/_0188_ ;
 wire \soc/spimemio/_0189_ ;
 wire \soc/spimemio/_0190_ ;
 wire \soc/spimemio/_0191_ ;
 wire \soc/spimemio/_0192_ ;
 wire \soc/spimemio/_0193_ ;
 wire net295;
 wire \soc/spimemio/_0195_ ;
 wire \soc/spimemio/_0196_ ;
 wire \soc/spimemio/_0197_ ;
 wire \soc/spimemio/_0198_ ;
 wire \soc/spimemio/_0199_ ;
 wire \soc/spimemio/_0200_ ;
 wire \soc/spimemio/_0201_ ;
 wire \soc/spimemio/_0202_ ;
 wire \soc/spimemio/_0203_ ;
 wire \soc/spimemio/_0204_ ;
 wire \soc/spimemio/_0205_ ;
 wire \soc/spimemio/_0206_ ;
 wire \soc/spimemio/_0207_ ;
 wire \soc/spimemio/_0208_ ;
 wire \soc/spimemio/_0209_ ;
 wire \soc/spimemio/_0210_ ;
 wire \soc/spimemio/_0211_ ;
 wire \soc/spimemio/_0212_ ;
 wire \soc/spimemio/_0213_ ;
 wire \soc/spimemio/_0214_ ;
 wire \soc/spimemio/_0215_ ;
 wire \soc/spimemio/_0216_ ;
 wire \soc/spimemio/_0217_ ;
 wire \soc/spimemio/_0218_ ;
 wire \soc/spimemio/_0219_ ;
 wire \soc/spimemio/_0220_ ;
 wire \soc/spimemio/_0221_ ;
 wire \soc/spimemio/_0222_ ;
 wire \soc/spimemio/_0223_ ;
 wire \soc/spimemio/_0224_ ;
 wire \soc/spimemio/_0225_ ;
 wire \soc/spimemio/_0226_ ;
 wire \soc/spimemio/_0227_ ;
 wire \soc/spimemio/_0228_ ;
 wire \soc/spimemio/_0229_ ;
 wire \soc/spimemio/_0230_ ;
 wire \soc/spimemio/_0231_ ;
 wire \soc/spimemio/_0232_ ;
 wire \soc/spimemio/_0233_ ;
 wire \soc/spimemio/_0234_ ;
 wire \soc/spimemio/_0235_ ;
 wire \soc/spimemio/_0236_ ;
 wire \soc/spimemio/_0237_ ;
 wire \soc/spimemio/_0238_ ;
 wire \soc/spimemio/_0239_ ;
 wire \soc/spimemio/_0240_ ;
 wire \soc/spimemio/_0241_ ;
 wire \soc/spimemio/_0242_ ;
 wire \soc/spimemio/_0243_ ;
 wire \soc/spimemio/_0244_ ;
 wire \soc/spimemio/_0245_ ;
 wire \soc/spimemio/_0246_ ;
 wire net294;
 wire \soc/spimemio/_0248_ ;
 wire \soc/spimemio/_0249_ ;
 wire net293;
 wire \soc/spimemio/_0251_ ;
 wire \soc/spimemio/_0252_ ;
 wire net292;
 wire net291;
 wire \soc/spimemio/_0255_ ;
 wire net290;
 wire \soc/spimemio/_0257_ ;
 wire \soc/spimemio/_0258_ ;
 wire \soc/spimemio/_0259_ ;
 wire \soc/spimemio/_0260_ ;
 wire \soc/spimemio/_0261_ ;
 wire \soc/spimemio/_0262_ ;
 wire \soc/spimemio/_0263_ ;
 wire \soc/spimemio/_0264_ ;
 wire \soc/spimemio/_0265_ ;
 wire \soc/spimemio/_0266_ ;
 wire \soc/spimemio/_0267_ ;
 wire \soc/spimemio/_0268_ ;
 wire \soc/spimemio/_0269_ ;
 wire \soc/spimemio/_0270_ ;
 wire net289;
 wire \soc/spimemio/_0272_ ;
 wire \soc/spimemio/_0273_ ;
 wire \soc/spimemio/_0274_ ;
 wire net288;
 wire \soc/spimemio/_0276_ ;
 wire \soc/spimemio/_0277_ ;
 wire \soc/spimemio/_0278_ ;
 wire \soc/spimemio/_0279_ ;
 wire \soc/spimemio/_0280_ ;
 wire \soc/spimemio/_0281_ ;
 wire \soc/spimemio/_0282_ ;
 wire \soc/spimemio/_0283_ ;
 wire \soc/spimemio/_0284_ ;
 wire \soc/spimemio/_0285_ ;
 wire \soc/spimemio/_0286_ ;
 wire net287;
 wire net286;
 wire \soc/spimemio/_0289_ ;
 wire \soc/spimemio/_0290_ ;
 wire \soc/spimemio/_0291_ ;
 wire \soc/spimemio/_0292_ ;
 wire \soc/spimemio/_0293_ ;
 wire \soc/spimemio/_0294_ ;
 wire \soc/spimemio/_0295_ ;
 wire \soc/spimemio/_0296_ ;
 wire \soc/spimemio/_0297_ ;
 wire \soc/spimemio/_0298_ ;
 wire \soc/spimemio/_0299_ ;
 wire \soc/spimemio/_0300_ ;
 wire \soc/spimemio/_0301_ ;
 wire \soc/spimemio/_0302_ ;
 wire \soc/spimemio/_0303_ ;
 wire \soc/spimemio/_0304_ ;
 wire \soc/spimemio/_0305_ ;
 wire \soc/spimemio/_0306_ ;
 wire net285;
 wire \soc/spimemio/_0308_ ;
 wire \soc/spimemio/_0309_ ;
 wire net284;
 wire \soc/spimemio/_0311_ ;
 wire \soc/spimemio/_0312_ ;
 wire \soc/spimemio/_0313_ ;
 wire net283;
 wire \soc/spimemio/_0315_ ;
 wire \soc/spimemio/_0316_ ;
 wire \soc/spimemio/_0317_ ;
 wire net282;
 wire \soc/spimemio/_0319_ ;
 wire \soc/spimemio/_0320_ ;
 wire \soc/spimemio/_0321_ ;
 wire \soc/spimemio/_0322_ ;
 wire \soc/spimemio/_0323_ ;
 wire net281;
 wire \soc/spimemio/_0325_ ;
 wire \soc/spimemio/_0326_ ;
 wire \soc/spimemio/_0327_ ;
 wire \soc/spimemio/_0328_ ;
 wire net280;
 wire \soc/spimemio/_0330_ ;
 wire \soc/spimemio/_0331_ ;
 wire \soc/spimemio/_0332_ ;
 wire \soc/spimemio/_0333_ ;
 wire \soc/spimemio/_0334_ ;
 wire \soc/spimemio/_0335_ ;
 wire \soc/spimemio/_0336_ ;
 wire \soc/spimemio/_0337_ ;
 wire \soc/spimemio/_0338_ ;
 wire \soc/spimemio/_0339_ ;
 wire \soc/spimemio/_0340_ ;
 wire \soc/spimemio/_0341_ ;
 wire \soc/spimemio/_0342_ ;
 wire \soc/spimemio/_0343_ ;
 wire \soc/spimemio/_0344_ ;
 wire \soc/spimemio/_0345_ ;
 wire \soc/spimemio/_0346_ ;
 wire \soc/spimemio/_0347_ ;
 wire \soc/spimemio/_0348_ ;
 wire \soc/spimemio/_0349_ ;
 wire \soc/spimemio/_0350_ ;
 wire \soc/spimemio/_0351_ ;
 wire \soc/spimemio/_0352_ ;
 wire \soc/spimemio/_0353_ ;
 wire \soc/spimemio/_0354_ ;
 wire \soc/spimemio/_0355_ ;
 wire \soc/spimemio/_0356_ ;
 wire \soc/spimemio/_0357_ ;
 wire \soc/spimemio/_0358_ ;
 wire \soc/spimemio/_0359_ ;
 wire \soc/spimemio/_0360_ ;
 wire \soc/spimemio/_0361_ ;
 wire \soc/spimemio/_0362_ ;
 wire \soc/spimemio/_0363_ ;
 wire \soc/spimemio/_0364_ ;
 wire \soc/spimemio/_0365_ ;
 wire \soc/spimemio/_0366_ ;
 wire \soc/spimemio/_0367_ ;
 wire \soc/spimemio/_0368_ ;
 wire net279;
 wire net278;
 wire \soc/spimemio/_0371_ ;
 wire net277;
 wire \soc/spimemio/_0373_ ;
 wire \soc/spimemio/_0374_ ;
 wire \soc/spimemio/_0375_ ;
 wire \soc/spimemio/_0376_ ;
 wire \soc/spimemio/_0377_ ;
 wire \soc/spimemio/_0378_ ;
 wire \soc/spimemio/_0379_ ;
 wire \soc/spimemio/_0380_ ;
 wire \soc/spimemio/_0381_ ;
 wire \soc/spimemio/_0382_ ;
 wire \soc/spimemio/_0383_ ;
 wire \soc/spimemio/_0384_ ;
 wire \soc/spimemio/_0385_ ;
 wire \soc/spimemio/_0386_ ;
 wire \soc/spimemio/_0387_ ;
 wire \soc/spimemio/_0388_ ;
 wire \soc/spimemio/_0389_ ;
 wire \soc/spimemio/_0390_ ;
 wire \soc/spimemio/_0391_ ;
 wire net276;
 wire \soc/spimemio/_0393_ ;
 wire net275;
 wire \soc/spimemio/_0395_ ;
 wire \soc/spimemio/_0396_ ;
 wire \soc/spimemio/_0397_ ;
 wire \soc/spimemio/_0398_ ;
 wire \soc/spimemio/_0399_ ;
 wire \soc/spimemio/_0400_ ;
 wire \soc/spimemio/_0401_ ;
 wire \soc/spimemio/_0402_ ;
 wire \soc/spimemio/_0403_ ;
 wire \soc/spimemio/_0404_ ;
 wire \soc/spimemio/_0405_ ;
 wire \soc/spimemio/_0406_ ;
 wire \soc/spimemio/_0407_ ;
 wire \soc/spimemio/_0408_ ;
 wire \soc/spimemio/_0409_ ;
 wire \soc/spimemio/_0410_ ;
 wire \soc/spimemio/_0411_ ;
 wire \soc/spimemio/_0412_ ;
 wire \soc/spimemio/_0413_ ;
 wire net274;
 wire \soc/spimemio/_0415_ ;
 wire net273;
 wire \soc/spimemio/_0417_ ;
 wire \soc/spimemio/_0418_ ;
 wire \soc/spimemio/_0419_ ;
 wire \soc/spimemio/_0420_ ;
 wire \soc/spimemio/_0421_ ;
 wire \soc/spimemio/_0422_ ;
 wire \soc/spimemio/_0423_ ;
 wire \soc/spimemio/_0424_ ;
 wire \soc/spimemio/_0425_ ;
 wire \soc/spimemio/_0426_ ;
 wire \soc/spimemio/_0427_ ;
 wire \soc/spimemio/_0428_ ;
 wire \soc/spimemio/_0429_ ;
 wire \soc/spimemio/_0430_ ;
 wire \soc/spimemio/_0431_ ;
 wire \soc/spimemio/_0432_ ;
 wire \soc/spimemio/_0433_ ;
 wire \soc/spimemio/_0434_ ;
 wire \soc/spimemio/_0435_ ;
 wire \soc/spimemio/_0436_ ;
 wire \soc/spimemio/_0437_ ;
 wire \soc/spimemio/_0438_ ;
 wire \soc/spimemio/_0439_ ;
 wire \soc/spimemio/_0440_ ;
 wire \soc/spimemio/_0441_ ;
 wire \soc/spimemio/_0442_ ;
 wire \soc/spimemio/_0443_ ;
 wire \soc/spimemio/_0444_ ;
 wire \soc/spimemio/_0445_ ;
 wire \soc/spimemio/_0446_ ;
 wire \soc/spimemio/_0447_ ;
 wire \soc/spimemio/_0448_ ;
 wire net272;
 wire \soc/spimemio/_0450_ ;
 wire \soc/spimemio/_0451_ ;
 wire \soc/spimemio/_0452_ ;
 wire \soc/spimemio/_0453_ ;
 wire \soc/spimemio/_0454_ ;
 wire \soc/spimemio/_0455_ ;
 wire \soc/spimemio/_0456_ ;
 wire \soc/spimemio/_0457_ ;
 wire \soc/spimemio/_0458_ ;
 wire \soc/spimemio/_0459_ ;
 wire \soc/spimemio/_0460_ ;
 wire \soc/spimemio/_0461_ ;
 wire \soc/spimemio/_0462_ ;
 wire \soc/spimemio/_0463_ ;
 wire \soc/spimemio/_0464_ ;
 wire \soc/spimemio/_0465_ ;
 wire \soc/spimemio/_0466_ ;
 wire \soc/spimemio/_0467_ ;
 wire \soc/spimemio/_0468_ ;
 wire \soc/spimemio/_0469_ ;
 wire \soc/spimemio/_0470_ ;
 wire \soc/spimemio/_0471_ ;
 wire \soc/spimemio/_0472_ ;
 wire \soc/spimemio/_0473_ ;
 wire \soc/spimemio/_0474_ ;
 wire \soc/spimemio/_0475_ ;
 wire \soc/spimemio/_0476_ ;
 wire \soc/spimemio/_0477_ ;
 wire \soc/spimemio/_0478_ ;
 wire \soc/spimemio/_0479_ ;
 wire \soc/spimemio/_0480_ ;
 wire \soc/spimemio/_0481_ ;
 wire \soc/spimemio/_0482_ ;
 wire \soc/spimemio/_0483_ ;
 wire \soc/spimemio/_0484_ ;
 wire \soc/spimemio/_0485_ ;
 wire \soc/spimemio/_0486_ ;
 wire \soc/spimemio/_0487_ ;
 wire \soc/spimemio/_0488_ ;
 wire \soc/spimemio/_0489_ ;
 wire \soc/spimemio/_0490_ ;
 wire \soc/spimemio/_0491_ ;
 wire \soc/spimemio/_0492_ ;
 wire \soc/spimemio/_0493_ ;
 wire \soc/spimemio/_0494_ ;
 wire \soc/spimemio/_0495_ ;
 wire \soc/spimemio/_0496_ ;
 wire \soc/spimemio/_0497_ ;
 wire \soc/spimemio/_0498_ ;
 wire \soc/spimemio/_0499_ ;
 wire \soc/spimemio/_0500_ ;
 wire \soc/spimemio/_0501_ ;
 wire \soc/spimemio/_0502_ ;
 wire \soc/spimemio/_0503_ ;
 wire \soc/spimemio/_0504_ ;
 wire \soc/spimemio/_0505_ ;
 wire \soc/spimemio/_0506_ ;
 wire net271;
 wire net270;
 wire \soc/spimemio/_0509_ ;
 wire \soc/spimemio/_0510_ ;
 wire \soc/spimemio/_0511_ ;
 wire \soc/spimemio/_0512_ ;
 wire \soc/spimemio/_0513_ ;
 wire \soc/spimemio/_0514_ ;
 wire \soc/spimemio/_0515_ ;
 wire \soc/spimemio/_0516_ ;
 wire \soc/spimemio/_0517_ ;
 wire \soc/spimemio/_0518_ ;
 wire \soc/spimemio/_0519_ ;
 wire \soc/spimemio/_0520_ ;
 wire \soc/spimemio/_0521_ ;
 wire \soc/spimemio/_0522_ ;
 wire \soc/spimemio/_0523_ ;
 wire \soc/spimemio/_0524_ ;
 wire \soc/spimemio/_0525_ ;
 wire \soc/spimemio/_0526_ ;
 wire \soc/spimemio/_0527_ ;
 wire \soc/spimemio/_0528_ ;
 wire \soc/spimemio/_0529_ ;
 wire \soc/spimemio/_0530_ ;
 wire \soc/spimemio/_0531_ ;
 wire \soc/spimemio/_0532_ ;
 wire \soc/spimemio/_0533_ ;
 wire \soc/spimemio/_0534_ ;
 wire \soc/spimemio/_0535_ ;
 wire \soc/spimemio/_0536_ ;
 wire \soc/spimemio/_0537_ ;
 wire \soc/spimemio/_0538_ ;
 wire \soc/spimemio/_0539_ ;
 wire \soc/spimemio/_0540_ ;
 wire \soc/spimemio/_0541_ ;
 wire \soc/spimemio/_0542_ ;
 wire \soc/spimemio/_0543_ ;
 wire \soc/spimemio/_0544_ ;
 wire \soc/spimemio/_0545_ ;
 wire \soc/spimemio/_0546_ ;
 wire net474;
 wire \soc/spimemio/buffer[0] ;
 wire \soc/spimemio/buffer[10] ;
 wire \soc/spimemio/buffer[11] ;
 wire \soc/spimemio/buffer[12] ;
 wire \soc/spimemio/buffer[13] ;
 wire \soc/spimemio/buffer[14] ;
 wire \soc/spimemio/buffer[15] ;
 wire \soc/spimemio/buffer[16] ;
 wire \soc/spimemio/buffer[17] ;
 wire \soc/spimemio/buffer[18] ;
 wire \soc/spimemio/buffer[19] ;
 wire \soc/spimemio/buffer[1] ;
 wire \soc/spimemio/buffer[20] ;
 wire \soc/spimemio/buffer[21] ;
 wire \soc/spimemio/buffer[22] ;
 wire \soc/spimemio/buffer[23] ;
 wire \soc/spimemio/buffer[2] ;
 wire \soc/spimemio/buffer[3] ;
 wire \soc/spimemio/buffer[4] ;
 wire \soc/spimemio/buffer[5] ;
 wire \soc/spimemio/buffer[6] ;
 wire \soc/spimemio/buffer[7] ;
 wire \soc/spimemio/buffer[8] ;
 wire \soc/spimemio/buffer[9] ;
 wire \soc/spimemio/config_clk ;
 wire \soc/spimemio/config_cont ;
 wire \soc/spimemio/config_csb ;
 wire \soc/spimemio/config_ddr ;
 wire \soc/spimemio/config_do[0] ;
 wire \soc/spimemio/config_do[1] ;
 wire \soc/spimemio/config_do[2] ;
 wire \soc/spimemio/config_do[3] ;
 wire \soc/spimemio/config_en ;
 wire \soc/spimemio/config_oe[0] ;
 wire \soc/spimemio/config_oe[1] ;
 wire \soc/spimemio/config_oe[2] ;
 wire \soc/spimemio/config_oe[3] ;
 wire \soc/spimemio/config_qspi ;
 wire \soc/spimemio/din_data[0] ;
 wire \soc/spimemio/din_data[1] ;
 wire \soc/spimemio/din_data[2] ;
 wire \soc/spimemio/din_data[3] ;
 wire \soc/spimemio/din_data[4] ;
 wire \soc/spimemio/din_data[5] ;
 wire \soc/spimemio/din_data[6] ;
 wire \soc/spimemio/din_data[7] ;
 wire \soc/spimemio/din_ddr ;
 wire \soc/spimemio/din_qspi ;
 wire \soc/spimemio/din_rd ;
 wire net239;
 wire \soc/spimemio/din_tag[0] ;
 wire \soc/spimemio/din_tag[1] ;
 wire \soc/spimemio/din_tag[2] ;
 wire \soc/spimemio/din_valid ;
 wire \soc/spimemio/dout_data[0] ;
 wire \soc/spimemio/dout_data[1] ;
 wire \soc/spimemio/dout_data[2] ;
 wire \soc/spimemio/dout_data[3] ;
 wire \soc/spimemio/dout_data[4] ;
 wire \soc/spimemio/dout_data[5] ;
 wire \soc/spimemio/dout_data[6] ;
 wire \soc/spimemio/dout_data[7] ;
 wire \soc/spimemio/dout_tag[0] ;
 wire \soc/spimemio/dout_tag[1] ;
 wire \soc/spimemio/dout_tag[2] ;
 wire \soc/spimemio/dout_tag[3] ;
 wire \soc/spimemio/dout_valid ;
 wire \soc/spimemio/rd_addr[0] ;
 wire \soc/spimemio/rd_addr[10] ;
 wire \soc/spimemio/rd_addr[11] ;
 wire \soc/spimemio/rd_addr[12] ;
 wire \soc/spimemio/rd_addr[13] ;
 wire \soc/spimemio/rd_addr[14] ;
 wire \soc/spimemio/rd_addr[15] ;
 wire \soc/spimemio/rd_addr[16] ;
 wire \soc/spimemio/rd_addr[17] ;
 wire \soc/spimemio/rd_addr[18] ;
 wire \soc/spimemio/rd_addr[19] ;
 wire \soc/spimemio/rd_addr[1] ;
 wire \soc/spimemio/rd_addr[20] ;
 wire \soc/spimemio/rd_addr[21] ;
 wire \soc/spimemio/rd_addr[22] ;
 wire \soc/spimemio/rd_addr[23] ;
 wire \soc/spimemio/rd_addr[2] ;
 wire \soc/spimemio/rd_addr[3] ;
 wire \soc/spimemio/rd_addr[4] ;
 wire \soc/spimemio/rd_addr[5] ;
 wire \soc/spimemio/rd_addr[6] ;
 wire \soc/spimemio/rd_addr[7] ;
 wire \soc/spimemio/rd_addr[8] ;
 wire \soc/spimemio/rd_addr[9] ;
 wire \soc/spimemio/rd_inc ;
 wire \soc/spimemio/rd_valid ;
 wire \soc/spimemio/rd_wait ;
 wire \soc/spimemio/softreset ;
 wire \soc/spimemio/state[0] ;
 wire \soc/spimemio/state[10] ;
 wire \soc/spimemio/state[11] ;
 wire \soc/spimemio/state[12] ;
 wire \soc/spimemio/state[1] ;
 wire \soc/spimemio/state[2] ;
 wire \soc/spimemio/state[3] ;
 wire \soc/spimemio/state[4] ;
 wire \soc/spimemio/state[5] ;
 wire \soc/spimemio/state[6] ;
 wire \soc/spimemio/state[7] ;
 wire \soc/spimemio/state[8] ;
 wire \soc/spimemio/state[9] ;
 wire \soc/spimemio/xfer_clk ;
 wire \soc/spimemio/xfer_csb ;
 wire \soc/spimemio/xfer_ddr ;
 wire \soc/spimemio/xfer_dspi ;
 wire \soc/spimemio/xfer_io0_90 ;
 wire \soc/spimemio/xfer_io0_do ;
 wire \soc/spimemio/xfer_io0_oe ;
 wire \soc/spimemio/xfer_io1_90 ;
 wire \soc/spimemio/xfer_io1_do ;
 wire \soc/spimemio/xfer_io1_oe ;
 wire \soc/spimemio/xfer_io2_90 ;
 wire \soc/spimemio/xfer_io2_do ;
 wire \soc/spimemio/xfer_io2_oe ;
 wire \soc/spimemio/xfer_io3_90 ;
 wire \soc/spimemio/xfer_io3_do ;
 wire net230;
 wire \soc/spimemio/xfer_resetn ;
 wire \soc/spimemio/xfer/_000_ ;
 wire \soc/spimemio/xfer/_001_ ;
 wire \soc/spimemio/xfer/_002_ ;
 wire \soc/spimemio/xfer/_003_ ;
 wire \soc/spimemio/xfer/_004_ ;
 wire \soc/spimemio/xfer/_005_ ;
 wire \soc/spimemio/xfer/_006_ ;
 wire \soc/spimemio/xfer/_007_ ;
 wire \soc/spimemio/xfer/_008_ ;
 wire \soc/spimemio/xfer/_009_ ;
 wire \soc/spimemio/xfer/_010_ ;
 wire \soc/spimemio/xfer/_011_ ;
 wire \soc/spimemio/xfer/_012_ ;
 wire \soc/spimemio/xfer/_013_ ;
 wire \soc/spimemio/xfer/_014_ ;
 wire \soc/spimemio/xfer/_015_ ;
 wire \soc/spimemio/xfer/_016_ ;
 wire \soc/spimemio/xfer/_017_ ;
 wire \soc/spimemio/xfer/_018_ ;
 wire \soc/spimemio/xfer/_019_ ;
 wire \soc/spimemio/xfer/_020_ ;
 wire \soc/spimemio/xfer/_021_ ;
 wire \soc/spimemio/xfer/_022_ ;
 wire \soc/spimemio/xfer/_023_ ;
 wire \soc/spimemio/xfer/_024_ ;
 wire \soc/spimemio/xfer/_025_ ;
 wire \soc/spimemio/xfer/_026_ ;
 wire \soc/spimemio/xfer/_027_ ;
 wire \soc/spimemio/xfer/_028_ ;
 wire \soc/spimemio/xfer/_029_ ;
 wire \soc/spimemio/xfer/_030_ ;
 wire \soc/spimemio/xfer/_031_ ;
 wire \soc/spimemio/xfer/_032_ ;
 wire \soc/spimemio/xfer/_033_ ;
 wire \soc/spimemio/xfer/_034_ ;
 wire \soc/spimemio/xfer/_035_ ;
 wire \soc/spimemio/xfer/_036_ ;
 wire \soc/spimemio/xfer/_037_ ;
 wire \soc/spimemio/xfer/_038_ ;
 wire \soc/spimemio/xfer/_039_ ;
 wire \soc/spimemio/xfer/_040_ ;
 wire \soc/spimemio/xfer/_041_ ;
 wire \soc/spimemio/xfer/_042_ ;
 wire net241;
 wire \soc/spimemio/xfer/_044_ ;
 wire \soc/spimemio/xfer/_045_ ;
 wire net240;
 wire \soc/spimemio/xfer/_047_ ;
 wire \soc/spimemio/xfer/_048_ ;
 wire \soc/spimemio/xfer/_049_ ;
 wire \soc/spimemio/xfer/_050_ ;
 wire \soc/spimemio/xfer/_051_ ;
 wire net238;
 wire net237;
 wire \soc/spimemio/xfer/_054_ ;
 wire \soc/spimemio/xfer/_055_ ;
 wire \soc/spimemio/xfer/_056_ ;
 wire \soc/spimemio/xfer/_057_ ;
 wire net236;
 wire \soc/spimemio/xfer/_059_ ;
 wire \soc/spimemio/xfer/_060_ ;
 wire \soc/spimemio/xfer/_061_ ;
 wire net235;
 wire \soc/spimemio/xfer/_063_ ;
 wire \soc/spimemio/xfer/_064_ ;
 wire \soc/spimemio/xfer/_065_ ;
 wire net234;
 wire net233;
 wire \soc/spimemio/xfer/_068_ ;
 wire \soc/spimemio/xfer/_069_ ;
 wire \soc/spimemio/xfer/_070_ ;
 wire \soc/spimemio/xfer/_071_ ;
 wire net232;
 wire \soc/spimemio/xfer/_073_ ;
 wire \soc/spimemio/xfer/_074_ ;
 wire \soc/spimemio/xfer/_075_ ;
 wire \soc/spimemio/xfer/_076_ ;
 wire \soc/spimemio/xfer/_077_ ;
 wire \soc/spimemio/xfer/_078_ ;
 wire \soc/spimemio/xfer/_079_ ;
 wire net231;
 wire \soc/spimemio/xfer/_081_ ;
 wire \soc/spimemio/xfer/_082_ ;
 wire \soc/spimemio/xfer/_083_ ;
 wire \soc/spimemio/xfer/_084_ ;
 wire \soc/spimemio/xfer/_085_ ;
 wire \soc/spimemio/xfer/_086_ ;
 wire \soc/spimemio/xfer/_087_ ;
 wire \soc/spimemio/xfer/_088_ ;
 wire \soc/spimemio/xfer/_089_ ;
 wire \soc/spimemio/xfer/_090_ ;
 wire \soc/spimemio/xfer/_091_ ;
 wire \soc/spimemio/xfer/_092_ ;
 wire \soc/spimemio/xfer/_093_ ;
 wire \soc/spimemio/xfer/_094_ ;
 wire \soc/spimemio/xfer/_095_ ;
 wire \soc/spimemio/xfer/_096_ ;
 wire \soc/spimemio/xfer/_097_ ;
 wire \soc/spimemio/xfer/_098_ ;
 wire \soc/spimemio/xfer/_099_ ;
 wire \soc/spimemio/xfer/_100_ ;
 wire \soc/spimemio/xfer/_101_ ;
 wire \soc/spimemio/xfer/_102_ ;
 wire \soc/spimemio/xfer/_103_ ;
 wire \soc/spimemio/xfer/_104_ ;
 wire \soc/spimemio/xfer/_105_ ;
 wire \soc/spimemio/xfer/_106_ ;
 wire \soc/spimemio/xfer/_107_ ;
 wire \soc/spimemio/xfer/_108_ ;
 wire \soc/spimemio/xfer/_109_ ;
 wire \soc/spimemio/xfer/_110_ ;
 wire \soc/spimemio/xfer/_111_ ;
 wire \soc/spimemio/xfer/_112_ ;
 wire \soc/spimemio/xfer/_113_ ;
 wire \soc/spimemio/xfer/_114_ ;
 wire \soc/spimemio/xfer/_115_ ;
 wire \soc/spimemio/xfer/_116_ ;
 wire \soc/spimemio/xfer/_117_ ;
 wire \soc/spimemio/xfer/_118_ ;
 wire \soc/spimemio/xfer/_119_ ;
 wire \soc/spimemio/xfer/_120_ ;
 wire \soc/spimemio/xfer/_121_ ;
 wire \soc/spimemio/xfer/_122_ ;
 wire \soc/spimemio/xfer/_123_ ;
 wire \soc/spimemio/xfer/_124_ ;
 wire \soc/spimemio/xfer/_125_ ;
 wire \soc/spimemio/xfer/_126_ ;
 wire \soc/spimemio/xfer/_127_ ;
 wire \soc/spimemio/xfer/_128_ ;
 wire \soc/spimemio/xfer/_129_ ;
 wire \soc/spimemio/xfer/_130_ ;
 wire \soc/spimemio/xfer/_131_ ;
 wire \soc/spimemio/xfer/_132_ ;
 wire \soc/spimemio/xfer/_133_ ;
 wire \soc/spimemio/xfer/_134_ ;
 wire \soc/spimemio/xfer/_135_ ;
 wire \soc/spimemio/xfer/_136_ ;
 wire \soc/spimemio/xfer/_137_ ;
 wire \soc/spimemio/xfer/_138_ ;
 wire \soc/spimemio/xfer/_139_ ;
 wire \soc/spimemio/xfer/_140_ ;
 wire \soc/spimemio/xfer/_141_ ;
 wire \soc/spimemio/xfer/_142_ ;
 wire \soc/spimemio/xfer/_143_ ;
 wire \soc/spimemio/xfer/_144_ ;
 wire \soc/spimemio/xfer/_145_ ;
 wire \soc/spimemio/xfer/_146_ ;
 wire \soc/spimemio/xfer/_147_ ;
 wire \soc/spimemio/xfer/_148_ ;
 wire \soc/spimemio/xfer/_149_ ;
 wire \soc/spimemio/xfer/_150_ ;
 wire \soc/spimemio/xfer/_151_ ;
 wire \soc/spimemio/xfer/_152_ ;
 wire \soc/spimemio/xfer/_153_ ;
 wire \soc/spimemio/xfer/_154_ ;
 wire \soc/spimemio/xfer/_155_ ;
 wire \soc/spimemio/xfer/_156_ ;
 wire \soc/spimemio/xfer/_157_ ;
 wire \soc/spimemio/xfer/_158_ ;
 wire \soc/spimemio/xfer/_159_ ;
 wire \soc/spimemio/xfer/_160_ ;
 wire \soc/spimemio/xfer/_161_ ;
 wire \soc/spimemio/xfer/_162_ ;
 wire \soc/spimemio/xfer/_163_ ;
 wire \soc/spimemio/xfer/_164_ ;
 wire \soc/spimemio/xfer/_165_ ;
 wire \soc/spimemio/xfer/_166_ ;
 wire \soc/spimemio/xfer/_167_ ;
 wire \soc/spimemio/xfer/_168_ ;
 wire \soc/spimemio/xfer/_169_ ;
 wire \soc/spimemio/xfer/_170_ ;
 wire \soc/spimemio/xfer/_171_ ;
 wire \soc/spimemio/xfer/_172_ ;
 wire \soc/spimemio/xfer/_173_ ;
 wire \soc/spimemio/xfer/_174_ ;
 wire \soc/spimemio/xfer/_175_ ;
 wire \soc/spimemio/xfer/_176_ ;
 wire \soc/spimemio/xfer/_177_ ;
 wire \soc/spimemio/xfer/_178_ ;
 wire \soc/spimemio/xfer/count[0] ;
 wire \soc/spimemio/xfer/count[1] ;
 wire \soc/spimemio/xfer/count[2] ;
 wire \soc/spimemio/xfer/count[3] ;
 wire \soc/spimemio/xfer/dummy_count[0] ;
 wire \soc/spimemio/xfer/dummy_count[1] ;
 wire \soc/spimemio/xfer/dummy_count[2] ;
 wire \soc/spimemio/xfer/dummy_count[3] ;
 wire \soc/spimemio/xfer/fetch ;
 wire \soc/spimemio/xfer/last_fetch ;
 wire \soc/spimemio/xfer/obuffer[0] ;
 wire \soc/spimemio/xfer/obuffer[1] ;
 wire \soc/spimemio/xfer/obuffer[2] ;
 wire \soc/spimemio/xfer/obuffer[3] ;
 wire \soc/spimemio/xfer/obuffer[4] ;
 wire \soc/spimemio/xfer/obuffer[5] ;
 wire \soc/spimemio/xfer/obuffer[6] ;
 wire \soc/spimemio/xfer/obuffer[7] ;
 wire \soc/spimemio/xfer/xfer_ddr ;
 wire \soc/spimemio/xfer/xfer_ddr_q ;
 wire \soc/spimemio/xfer/xfer_dspi ;
 wire \soc/spimemio/xfer/xfer_qspi ;
 wire \soc/spimemio/xfer/xfer_rd ;
 wire \soc/spimemio/xfer/xfer_tag[0] ;
 wire \soc/spimemio/xfer/xfer_tag[1] ;
 wire \soc/spimemio/xfer/xfer_tag[2] ;
 wire \soc/spimemio/xfer/xfer_tag[3] ;
 wire \wave_gen_inst/_0000_ ;
 wire \wave_gen_inst/_0001_ ;
 wire \wave_gen_inst/_0002_ ;
 wire \wave_gen_inst/_0003_ ;
 wire \wave_gen_inst/_0004_ ;
 wire \wave_gen_inst/_0005_ ;
 wire \wave_gen_inst/_0006_ ;
 wire \wave_gen_inst/_0007_ ;
 wire \wave_gen_inst/_0008_ ;
 wire \wave_gen_inst/_0009_ ;
 wire \wave_gen_inst/_0010_ ;
 wire \wave_gen_inst/_0011_ ;
 wire \wave_gen_inst/_0012_ ;
 wire \wave_gen_inst/_0013_ ;
 wire \wave_gen_inst/_0014_ ;
 wire \wave_gen_inst/_0015_ ;
 wire \wave_gen_inst/_0016_ ;
 wire \wave_gen_inst/_0017_ ;
 wire \wave_gen_inst/_0018_ ;
 wire \wave_gen_inst/_0019_ ;
 wire \wave_gen_inst/_0020_ ;
 wire \wave_gen_inst/_0021_ ;
 wire \wave_gen_inst/_0022_ ;
 wire \wave_gen_inst/_0023_ ;
 wire \wave_gen_inst/_0024_ ;
 wire \wave_gen_inst/_0025_ ;
 wire \wave_gen_inst/_0026_ ;
 wire \wave_gen_inst/_0027_ ;
 wire \wave_gen_inst/_0028_ ;
 wire \wave_gen_inst/_0029_ ;
 wire \wave_gen_inst/_0030_ ;
 wire \wave_gen_inst/_0031_ ;
 wire \wave_gen_inst/_0032_ ;
 wire \wave_gen_inst/_0033_ ;
 wire \wave_gen_inst/_0034_ ;
 wire \wave_gen_inst/_0035_ ;
 wire \wave_gen_inst/_0036_ ;
 wire \wave_gen_inst/_0037_ ;
 wire \wave_gen_inst/_0038_ ;
 wire \wave_gen_inst/_0039_ ;
 wire \wave_gen_inst/_0040_ ;
 wire \wave_gen_inst/_0041_ ;
 wire \wave_gen_inst/_0042_ ;
 wire \wave_gen_inst/_0043_ ;
 wire \wave_gen_inst/_0044_ ;
 wire \wave_gen_inst/_0045_ ;
 wire \wave_gen_inst/_0046_ ;
 wire \wave_gen_inst/_0047_ ;
 wire \wave_gen_inst/_0048_ ;
 wire \wave_gen_inst/_0049_ ;
 wire \wave_gen_inst/_0050_ ;
 wire \wave_gen_inst/_0051_ ;
 wire \wave_gen_inst/_0052_ ;
 wire \wave_gen_inst/_0053_ ;
 wire \wave_gen_inst/_0054_ ;
 wire \wave_gen_inst/_0055_ ;
 wire \wave_gen_inst/_0056_ ;
 wire \wave_gen_inst/_0057_ ;
 wire \wave_gen_inst/_0058_ ;
 wire \wave_gen_inst/_0059_ ;
 wire \wave_gen_inst/_0060_ ;
 wire \wave_gen_inst/_0061_ ;
 wire \wave_gen_inst/_0062_ ;
 wire \wave_gen_inst/_0063_ ;
 wire \wave_gen_inst/_0064_ ;
 wire \wave_gen_inst/_0065_ ;
 wire \wave_gen_inst/_0066_ ;
 wire \wave_gen_inst/_0067_ ;
 wire \wave_gen_inst/_0068_ ;
 wire \wave_gen_inst/_0069_ ;
 wire \wave_gen_inst/_0070_ ;
 wire \wave_gen_inst/_0071_ ;
 wire \wave_gen_inst/_0072_ ;
 wire \wave_gen_inst/_0073_ ;
 wire \wave_gen_inst/_0074_ ;
 wire \wave_gen_inst/_0075_ ;
 wire \wave_gen_inst/_0076_ ;
 wire \wave_gen_inst/_0077_ ;
 wire \wave_gen_inst/_0078_ ;
 wire \wave_gen_inst/_0079_ ;
 wire \wave_gen_inst/_0080_ ;
 wire \wave_gen_inst/_0081_ ;
 wire \wave_gen_inst/_0082_ ;
 wire \wave_gen_inst/_0083_ ;
 wire \wave_gen_inst/_0084_ ;
 wire \wave_gen_inst/_0085_ ;
 wire \wave_gen_inst/_0086_ ;
 wire \wave_gen_inst/_0087_ ;
 wire \wave_gen_inst/_0088_ ;
 wire \wave_gen_inst/_0089_ ;
 wire \wave_gen_inst/_0090_ ;
 wire \wave_gen_inst/_0091_ ;
 wire \wave_gen_inst/_0092_ ;
 wire \wave_gen_inst/_0093_ ;
 wire \wave_gen_inst/_0094_ ;
 wire \wave_gen_inst/_0095_ ;
 wire \wave_gen_inst/_0096_ ;
 wire \wave_gen_inst/_0097_ ;
 wire \wave_gen_inst/_0098_ ;
 wire \wave_gen_inst/_0099_ ;
 wire \wave_gen_inst/_0100_ ;
 wire \wave_gen_inst/_0101_ ;
 wire \wave_gen_inst/_0102_ ;
 wire \wave_gen_inst/_0103_ ;
 wire \wave_gen_inst/_0104_ ;
 wire \wave_gen_inst/_0105_ ;
 wire \wave_gen_inst/_0106_ ;
 wire net111;
 wire \wave_gen_inst/_0108_ ;
 wire \wave_gen_inst/_0109_ ;
 wire \wave_gen_inst/_0110_ ;
 wire \wave_gen_inst/_0111_ ;
 wire \wave_gen_inst/_0112_ ;
 wire \wave_gen_inst/_0113_ ;
 wire \wave_gen_inst/_0114_ ;
 wire \wave_gen_inst/_0115_ ;
 wire \wave_gen_inst/_0116_ ;
 wire \wave_gen_inst/_0117_ ;
 wire \wave_gen_inst/_0118_ ;
 wire \wave_gen_inst/_0119_ ;
 wire \wave_gen_inst/_0120_ ;
 wire \wave_gen_inst/_0121_ ;
 wire \wave_gen_inst/_0122_ ;
 wire \wave_gen_inst/_0123_ ;
 wire \wave_gen_inst/_0124_ ;
 wire \wave_gen_inst/_0125_ ;
 wire \wave_gen_inst/_0126_ ;
 wire \wave_gen_inst/_0127_ ;
 wire \wave_gen_inst/_0128_ ;
 wire \wave_gen_inst/_0129_ ;
 wire \wave_gen_inst/_0130_ ;
 wire \wave_gen_inst/_0131_ ;
 wire \wave_gen_inst/_0132_ ;
 wire \wave_gen_inst/_0133_ ;
 wire \wave_gen_inst/_0134_ ;
 wire \wave_gen_inst/_0135_ ;
 wire \wave_gen_inst/_0136_ ;
 wire \wave_gen_inst/_0137_ ;
 wire \wave_gen_inst/_0138_ ;
 wire \wave_gen_inst/_0139_ ;
 wire \wave_gen_inst/_0140_ ;
 wire \wave_gen_inst/_0141_ ;
 wire \wave_gen_inst/_0142_ ;
 wire \wave_gen_inst/_0143_ ;
 wire \wave_gen_inst/_0144_ ;
 wire \wave_gen_inst/_0145_ ;
 wire \wave_gen_inst/_0146_ ;
 wire \wave_gen_inst/_0147_ ;
 wire \wave_gen_inst/_0148_ ;
 wire \wave_gen_inst/_0149_ ;
 wire net110;
 wire \wave_gen_inst/_0151_ ;
 wire \wave_gen_inst/_0152_ ;
 wire \wave_gen_inst/_0153_ ;
 wire \wave_gen_inst/_0154_ ;
 wire \wave_gen_inst/_0155_ ;
 wire \wave_gen_inst/_0156_ ;
 wire \wave_gen_inst/_0157_ ;
 wire net109;
 wire \wave_gen_inst/_0159_ ;
 wire \wave_gen_inst/_0160_ ;
 wire \wave_gen_inst/_0161_ ;
 wire \wave_gen_inst/_0162_ ;
 wire \wave_gen_inst/_0163_ ;
 wire \wave_gen_inst/_0164_ ;
 wire net108;
 wire \wave_gen_inst/_0166_ ;
 wire \wave_gen_inst/_0167_ ;
 wire net107;
 wire \wave_gen_inst/_0169_ ;
 wire net106;
 wire \wave_gen_inst/_0171_ ;
 wire net105;
 wire net104;
 wire \wave_gen_inst/_0174_ ;
 wire \wave_gen_inst/_0175_ ;
 wire \wave_gen_inst/_0176_ ;
 wire \wave_gen_inst/_0177_ ;
 wire \wave_gen_inst/_0178_ ;
 wire \wave_gen_inst/_0179_ ;
 wire \wave_gen_inst/_0180_ ;
 wire \wave_gen_inst/_0181_ ;
 wire \wave_gen_inst/_0182_ ;
 wire \wave_gen_inst/_0183_ ;
 wire \wave_gen_inst/_0184_ ;
 wire \wave_gen_inst/_0185_ ;
 wire \wave_gen_inst/_0186_ ;
 wire \wave_gen_inst/_0187_ ;
 wire \wave_gen_inst/_0188_ ;
 wire \wave_gen_inst/_0189_ ;
 wire \wave_gen_inst/_0190_ ;
 wire \wave_gen_inst/_0191_ ;
 wire \wave_gen_inst/_0192_ ;
 wire \wave_gen_inst/_0193_ ;
 wire \wave_gen_inst/_0194_ ;
 wire \wave_gen_inst/_0195_ ;
 wire \wave_gen_inst/_0196_ ;
 wire \wave_gen_inst/_0197_ ;
 wire \wave_gen_inst/_0198_ ;
 wire \wave_gen_inst/_0199_ ;
 wire \wave_gen_inst/_0200_ ;
 wire \wave_gen_inst/_0201_ ;
 wire \wave_gen_inst/_0202_ ;
 wire \wave_gen_inst/_0203_ ;
 wire \wave_gen_inst/_0204_ ;
 wire \wave_gen_inst/_0205_ ;
 wire \wave_gen_inst/_0206_ ;
 wire \wave_gen_inst/_0207_ ;
 wire \wave_gen_inst/_0208_ ;
 wire \wave_gen_inst/_0209_ ;
 wire \wave_gen_inst/_0210_ ;
 wire \wave_gen_inst/_0211_ ;
 wire \wave_gen_inst/_0212_ ;
 wire \wave_gen_inst/_0213_ ;
 wire \wave_gen_inst/_0214_ ;
 wire \wave_gen_inst/_0215_ ;
 wire \wave_gen_inst/_0216_ ;
 wire \wave_gen_inst/_0217_ ;
 wire \wave_gen_inst/_0218_ ;
 wire \wave_gen_inst/_0219_ ;
 wire \wave_gen_inst/_0220_ ;
 wire \wave_gen_inst/_0221_ ;
 wire \wave_gen_inst/_0222_ ;
 wire \wave_gen_inst/_0223_ ;
 wire \wave_gen_inst/_0224_ ;
 wire \wave_gen_inst/_0225_ ;
 wire \wave_gen_inst/_0226_ ;
 wire \wave_gen_inst/_0227_ ;
 wire \wave_gen_inst/_0228_ ;
 wire \wave_gen_inst/_0229_ ;
 wire \wave_gen_inst/_0230_ ;
 wire \wave_gen_inst/_0231_ ;
 wire \wave_gen_inst/_0232_ ;
 wire \wave_gen_inst/_0233_ ;
 wire \wave_gen_inst/_0234_ ;
 wire \wave_gen_inst/_0235_ ;
 wire \wave_gen_inst/_0236_ ;
 wire \wave_gen_inst/_0237_ ;
 wire \wave_gen_inst/_0238_ ;
 wire \wave_gen_inst/_0239_ ;
 wire \wave_gen_inst/_0240_ ;
 wire \wave_gen_inst/_0241_ ;
 wire \wave_gen_inst/_0242_ ;
 wire \wave_gen_inst/_0243_ ;
 wire \wave_gen_inst/_0244_ ;
 wire \wave_gen_inst/_0245_ ;
 wire \wave_gen_inst/_0246_ ;
 wire \wave_gen_inst/_0247_ ;
 wire \wave_gen_inst/_0248_ ;
 wire net103;
 wire \wave_gen_inst/_0250_ ;
 wire \wave_gen_inst/_0251_ ;
 wire \wave_gen_inst/_0252_ ;
 wire \wave_gen_inst/_0253_ ;
 wire \wave_gen_inst/_0254_ ;
 wire \wave_gen_inst/_0255_ ;
 wire \wave_gen_inst/_0256_ ;
 wire \wave_gen_inst/_0257_ ;
 wire \wave_gen_inst/_0258_ ;
 wire \wave_gen_inst/_0259_ ;
 wire \wave_gen_inst/_0260_ ;
 wire \wave_gen_inst/_0261_ ;
 wire \wave_gen_inst/_0262_ ;
 wire \wave_gen_inst/_0263_ ;
 wire \wave_gen_inst/_0264_ ;
 wire \wave_gen_inst/_0265_ ;
 wire \wave_gen_inst/_0266_ ;
 wire \wave_gen_inst/_0267_ ;
 wire \wave_gen_inst/_0268_ ;
 wire \wave_gen_inst/_0269_ ;
 wire \wave_gen_inst/_0270_ ;
 wire \wave_gen_inst/_0271_ ;
 wire \wave_gen_inst/_0272_ ;
 wire \wave_gen_inst/_0273_ ;
 wire \wave_gen_inst/_0274_ ;
 wire \wave_gen_inst/_0275_ ;
 wire net102;
 wire \wave_gen_inst/_0277_ ;
 wire \wave_gen_inst/_0278_ ;
 wire \wave_gen_inst/_0279_ ;
 wire \wave_gen_inst/_0280_ ;
 wire \wave_gen_inst/_0281_ ;
 wire \wave_gen_inst/_0282_ ;
 wire \wave_gen_inst/_0283_ ;
 wire \wave_gen_inst/_0284_ ;
 wire \wave_gen_inst/_0285_ ;
 wire \wave_gen_inst/_0286_ ;
 wire \wave_gen_inst/_0287_ ;
 wire \wave_gen_inst/_0288_ ;
 wire \wave_gen_inst/_0289_ ;
 wire \wave_gen_inst/_0290_ ;
 wire \wave_gen_inst/_0291_ ;
 wire \wave_gen_inst/_0292_ ;
 wire \wave_gen_inst/_0293_ ;
 wire \wave_gen_inst/_0294_ ;
 wire \wave_gen_inst/_0295_ ;
 wire \wave_gen_inst/_0296_ ;
 wire \wave_gen_inst/_0297_ ;
 wire \wave_gen_inst/_0298_ ;
 wire \wave_gen_inst/_0299_ ;
 wire \wave_gen_inst/_0300_ ;
 wire \wave_gen_inst/_0301_ ;
 wire \wave_gen_inst/_0302_ ;
 wire \wave_gen_inst/_0303_ ;
 wire \wave_gen_inst/_0304_ ;
 wire \wave_gen_inst/_0305_ ;
 wire \wave_gen_inst/_0306_ ;
 wire \wave_gen_inst/_0307_ ;
 wire \wave_gen_inst/_0308_ ;
 wire \wave_gen_inst/_0309_ ;
 wire \wave_gen_inst/_0310_ ;
 wire \wave_gen_inst/_0311_ ;
 wire \wave_gen_inst/_0312_ ;
 wire \wave_gen_inst/_0313_ ;
 wire \wave_gen_inst/_0314_ ;
 wire \wave_gen_inst/_0315_ ;
 wire \wave_gen_inst/_0316_ ;
 wire \wave_gen_inst/_0317_ ;
 wire \wave_gen_inst/_0318_ ;
 wire \wave_gen_inst/_0319_ ;
 wire \wave_gen_inst/_0320_ ;
 wire \wave_gen_inst/_0321_ ;
 wire \wave_gen_inst/_0322_ ;
 wire \wave_gen_inst/_0323_ ;
 wire \wave_gen_inst/_0324_ ;
 wire \wave_gen_inst/_0325_ ;
 wire \wave_gen_inst/_0326_ ;
 wire \wave_gen_inst/_0327_ ;
 wire \wave_gen_inst/_0328_ ;
 wire \wave_gen_inst/_0329_ ;
 wire \wave_gen_inst/_0330_ ;
 wire \wave_gen_inst/_0331_ ;
 wire \wave_gen_inst/_0332_ ;
 wire \wave_gen_inst/_0333_ ;
 wire \wave_gen_inst/_0334_ ;
 wire \wave_gen_inst/_0335_ ;
 wire \wave_gen_inst/_0336_ ;
 wire \wave_gen_inst/_0337_ ;
 wire \wave_gen_inst/_0338_ ;
 wire \wave_gen_inst/_0339_ ;
 wire \wave_gen_inst/_0340_ ;
 wire \wave_gen_inst/_0341_ ;
 wire \wave_gen_inst/_0342_ ;
 wire \wave_gen_inst/_0343_ ;
 wire \wave_gen_inst/_0344_ ;
 wire \wave_gen_inst/_0345_ ;
 wire \wave_gen_inst/_0346_ ;
 wire \wave_gen_inst/_0347_ ;
 wire \wave_gen_inst/_0348_ ;
 wire \wave_gen_inst/_0349_ ;
 wire \wave_gen_inst/_0350_ ;
 wire \wave_gen_inst/_0351_ ;
 wire \wave_gen_inst/_0352_ ;
 wire \wave_gen_inst/_0353_ ;
 wire \wave_gen_inst/_0354_ ;
 wire \wave_gen_inst/_0355_ ;
 wire \wave_gen_inst/_0356_ ;
 wire \wave_gen_inst/_0357_ ;
 wire \wave_gen_inst/_0358_ ;
 wire \wave_gen_inst/_0359_ ;
 wire \wave_gen_inst/_0360_ ;
 wire \wave_gen_inst/_0361_ ;
 wire \wave_gen_inst/_0362_ ;
 wire \wave_gen_inst/_0363_ ;
 wire \wave_gen_inst/_0364_ ;
 wire \wave_gen_inst/_0365_ ;
 wire \wave_gen_inst/_0366_ ;
 wire \wave_gen_inst/_0367_ ;
 wire \wave_gen_inst/_0368_ ;
 wire \wave_gen_inst/_0369_ ;
 wire \wave_gen_inst/_0370_ ;
 wire \wave_gen_inst/_0371_ ;
 wire \wave_gen_inst/_0372_ ;
 wire \wave_gen_inst/_0373_ ;
 wire net101;
 wire \wave_gen_inst/_0375_ ;
 wire \wave_gen_inst/_0376_ ;
 wire \wave_gen_inst/_0377_ ;
 wire \wave_gen_inst/_0378_ ;
 wire \wave_gen_inst/_0379_ ;
 wire \wave_gen_inst/_0380_ ;
 wire \wave_gen_inst/_0381_ ;
 wire \wave_gen_inst/_0382_ ;
 wire \wave_gen_inst/_0383_ ;
 wire \wave_gen_inst/_0384_ ;
 wire \wave_gen_inst/_0385_ ;
 wire \wave_gen_inst/_0386_ ;
 wire \wave_gen_inst/_0387_ ;
 wire \wave_gen_inst/_0388_ ;
 wire \wave_gen_inst/_0389_ ;
 wire \wave_gen_inst/_0390_ ;
 wire \wave_gen_inst/_0391_ ;
 wire \wave_gen_inst/_0392_ ;
 wire \wave_gen_inst/_0393_ ;
 wire \wave_gen_inst/_0394_ ;
 wire \wave_gen_inst/_0395_ ;
 wire \wave_gen_inst/_0396_ ;
 wire \wave_gen_inst/_0397_ ;
 wire \wave_gen_inst/_0398_ ;
 wire \wave_gen_inst/_0399_ ;
 wire \wave_gen_inst/_0400_ ;
 wire \wave_gen_inst/_0401_ ;
 wire \wave_gen_inst/_0402_ ;
 wire \wave_gen_inst/_0403_ ;
 wire \wave_gen_inst/_0404_ ;
 wire \wave_gen_inst/_0405_ ;
 wire \wave_gen_inst/_0406_ ;
 wire \wave_gen_inst/_0407_ ;
 wire \wave_gen_inst/_0408_ ;
 wire \wave_gen_inst/_0409_ ;
 wire \wave_gen_inst/_0410_ ;
 wire \wave_gen_inst/_0411_ ;
 wire \wave_gen_inst/_0412_ ;
 wire \wave_gen_inst/_0413_ ;
 wire \wave_gen_inst/_0414_ ;
 wire \wave_gen_inst/_0415_ ;
 wire \wave_gen_inst/_0416_ ;
 wire \wave_gen_inst/_0417_ ;
 wire \wave_gen_inst/_0418_ ;
 wire \wave_gen_inst/_0419_ ;
 wire \wave_gen_inst/_0420_ ;
 wire \wave_gen_inst/_0421_ ;
 wire \wave_gen_inst/_0422_ ;
 wire \wave_gen_inst/_0423_ ;
 wire \wave_gen_inst/_0424_ ;
 wire \wave_gen_inst/_0425_ ;
 wire \wave_gen_inst/_0426_ ;
 wire \wave_gen_inst/_0427_ ;
 wire \wave_gen_inst/_0428_ ;
 wire \wave_gen_inst/_0429_ ;
 wire \wave_gen_inst/_0430_ ;
 wire \wave_gen_inst/_0431_ ;
 wire \wave_gen_inst/_0432_ ;
 wire \wave_gen_inst/_0433_ ;
 wire \wave_gen_inst/_0434_ ;
 wire \wave_gen_inst/_0435_ ;
 wire \wave_gen_inst/_0436_ ;
 wire \wave_gen_inst/_0437_ ;
 wire \wave_gen_inst/_0438_ ;
 wire \wave_gen_inst/_0439_ ;
 wire \wave_gen_inst/_0440_ ;
 wire \wave_gen_inst/_0441_ ;
 wire \wave_gen_inst/_0442_ ;
 wire \wave_gen_inst/_0443_ ;
 wire \wave_gen_inst/_0444_ ;
 wire \wave_gen_inst/_0445_ ;
 wire \wave_gen_inst/_0446_ ;
 wire \wave_gen_inst/_0447_ ;
 wire \wave_gen_inst/_0448_ ;
 wire \wave_gen_inst/_0449_ ;
 wire \wave_gen_inst/_0450_ ;
 wire net100;
 wire net99;
 wire net98;
 wire \wave_gen_inst/_0454_ ;
 wire \wave_gen_inst/_0455_ ;
 wire \wave_gen_inst/_0456_ ;
 wire \wave_gen_inst/_0457_ ;
 wire \wave_gen_inst/_0458_ ;
 wire \wave_gen_inst/_0459_ ;
 wire \wave_gen_inst/_0460_ ;
 wire \wave_gen_inst/_0461_ ;
 wire \wave_gen_inst/_0462_ ;
 wire \wave_gen_inst/_0463_ ;
 wire \wave_gen_inst/_0464_ ;
 wire \wave_gen_inst/_0465_ ;
 wire \wave_gen_inst/_0466_ ;
 wire \wave_gen_inst/_0467_ ;
 wire \wave_gen_inst/_0468_ ;
 wire \wave_gen_inst/_0469_ ;
 wire \wave_gen_inst/_0470_ ;
 wire \wave_gen_inst/_0471_ ;
 wire \wave_gen_inst/_0472_ ;
 wire \wave_gen_inst/_0473_ ;
 wire \wave_gen_inst/_0474_ ;
 wire \wave_gen_inst/_0475_ ;
 wire \wave_gen_inst/_0476_ ;
 wire \wave_gen_inst/_0477_ ;
 wire \wave_gen_inst/_0478_ ;
 wire \wave_gen_inst/_0479_ ;
 wire \wave_gen_inst/_0480_ ;
 wire \wave_gen_inst/_0481_ ;
 wire \wave_gen_inst/_0482_ ;
 wire \wave_gen_inst/_0483_ ;
 wire \wave_gen_inst/_0484_ ;
 wire \wave_gen_inst/_0485_ ;
 wire \wave_gen_inst/_0486_ ;
 wire \wave_gen_inst/_0487_ ;
 wire \wave_gen_inst/_0488_ ;
 wire \wave_gen_inst/_0489_ ;
 wire \wave_gen_inst/_0490_ ;
 wire \wave_gen_inst/_0491_ ;
 wire \wave_gen_inst/_0492_ ;
 wire \wave_gen_inst/_0493_ ;
 wire \wave_gen_inst/_0494_ ;
 wire \wave_gen_inst/_0495_ ;
 wire \wave_gen_inst/_0496_ ;
 wire \wave_gen_inst/_0497_ ;
 wire \wave_gen_inst/_0498_ ;
 wire \wave_gen_inst/_0499_ ;
 wire \wave_gen_inst/_0500_ ;
 wire \wave_gen_inst/_0501_ ;
 wire \wave_gen_inst/_0502_ ;
 wire \wave_gen_inst/_0503_ ;
 wire \wave_gen_inst/_0504_ ;
 wire \wave_gen_inst/_0505_ ;
 wire \wave_gen_inst/_0506_ ;
 wire \wave_gen_inst/_0507_ ;
 wire \wave_gen_inst/_0508_ ;
 wire \wave_gen_inst/_0509_ ;
 wire \wave_gen_inst/_0510_ ;
 wire \wave_gen_inst/_0511_ ;
 wire \wave_gen_inst/_0512_ ;
 wire \wave_gen_inst/_0513_ ;
 wire \wave_gen_inst/_0514_ ;
 wire \wave_gen_inst/_0515_ ;
 wire \wave_gen_inst/_0516_ ;
 wire \wave_gen_inst/_0517_ ;
 wire \wave_gen_inst/_0518_ ;
 wire \wave_gen_inst/_0519_ ;
 wire \wave_gen_inst/_0520_ ;
 wire \wave_gen_inst/_0521_ ;
 wire \wave_gen_inst/_0522_ ;
 wire \wave_gen_inst/_0523_ ;
 wire \wave_gen_inst/_0524_ ;
 wire \wave_gen_inst/_0525_ ;
 wire \wave_gen_inst/_0526_ ;
 wire \wave_gen_inst/_0527_ ;
 wire \wave_gen_inst/_0528_ ;
 wire \wave_gen_inst/_0529_ ;
 wire \wave_gen_inst/_0530_ ;
 wire \wave_gen_inst/_0531_ ;
 wire \wave_gen_inst/_0532_ ;
 wire \wave_gen_inst/_0533_ ;
 wire \wave_gen_inst/_0534_ ;
 wire \wave_gen_inst/_0535_ ;
 wire \wave_gen_inst/_0536_ ;
 wire \wave_gen_inst/_0537_ ;
 wire \wave_gen_inst/_0538_ ;
 wire \wave_gen_inst/_0539_ ;
 wire \wave_gen_inst/_0540_ ;
 wire \wave_gen_inst/_0541_ ;
 wire \wave_gen_inst/_0542_ ;
 wire \wave_gen_inst/_0543_ ;
 wire \wave_gen_inst/_0544_ ;
 wire \wave_gen_inst/_0545_ ;
 wire \wave_gen_inst/_0546_ ;
 wire \wave_gen_inst/_0547_ ;
 wire \wave_gen_inst/_0548_ ;
 wire \wave_gen_inst/_0549_ ;
 wire \wave_gen_inst/_0550_ ;
 wire \wave_gen_inst/_0551_ ;
 wire \wave_gen_inst/_0552_ ;
 wire \wave_gen_inst/_0553_ ;
 wire \wave_gen_inst/_0554_ ;
 wire \wave_gen_inst/_0555_ ;
 wire \wave_gen_inst/_0556_ ;
 wire \wave_gen_inst/_0557_ ;
 wire \wave_gen_inst/_0558_ ;
 wire \wave_gen_inst/_0559_ ;
 wire \wave_gen_inst/_0560_ ;
 wire \wave_gen_inst/_0561_ ;
 wire \wave_gen_inst/_0562_ ;
 wire \wave_gen_inst/_0563_ ;
 wire \wave_gen_inst/_0564_ ;
 wire \wave_gen_inst/_0565_ ;
 wire \wave_gen_inst/_0566_ ;
 wire \wave_gen_inst/_0567_ ;
 wire net97;
 wire net96;
 wire \wave_gen_inst/_0570_ ;
 wire net95;
 wire net94;
 wire \wave_gen_inst/_0573_ ;
 wire \wave_gen_inst/_0574_ ;
 wire \wave_gen_inst/_0575_ ;
 wire \wave_gen_inst/_0576_ ;
 wire \wave_gen_inst/_0577_ ;
 wire \wave_gen_inst/_0578_ ;
 wire \wave_gen_inst/_0579_ ;
 wire \wave_gen_inst/_0580_ ;
 wire net93;
 wire \wave_gen_inst/_0582_ ;
 wire \wave_gen_inst/_0583_ ;
 wire \wave_gen_inst/_0584_ ;
 wire \wave_gen_inst/_0585_ ;
 wire net92;
 wire \wave_gen_inst/_0587_ ;
 wire net91;
 wire \wave_gen_inst/_0589_ ;
 wire net90;
 wire \wave_gen_inst/_0591_ ;
 wire net89;
 wire \wave_gen_inst/_0593_ ;
 wire net88;
 wire \wave_gen_inst/_0595_ ;
 wire net87;
 wire \wave_gen_inst/_0597_ ;
 wire net86;
 wire net85;
 wire \wave_gen_inst/_0600_ ;
 wire \wave_gen_inst/_0601_ ;
 wire \wave_gen_inst/_0602_ ;
 wire net84;
 wire net83;
 wire \wave_gen_inst/_0605_ ;
 wire \wave_gen_inst/_0606_ ;
 wire \wave_gen_inst/_0607_ ;
 wire \wave_gen_inst/_0608_ ;
 wire \wave_gen_inst/_0609_ ;
 wire \wave_gen_inst/_0610_ ;
 wire \wave_gen_inst/_0611_ ;
 wire \wave_gen_inst/_0612_ ;
 wire \wave_gen_inst/_0613_ ;
 wire \wave_gen_inst/_0614_ ;
 wire \wave_gen_inst/_0615_ ;
 wire \wave_gen_inst/_0616_ ;
 wire \wave_gen_inst/_0617_ ;
 wire \wave_gen_inst/_0618_ ;
 wire \wave_gen_inst/_0619_ ;
 wire \wave_gen_inst/_0620_ ;
 wire \wave_gen_inst/_0621_ ;
 wire \wave_gen_inst/_0622_ ;
 wire \wave_gen_inst/_0623_ ;
 wire \wave_gen_inst/_0624_ ;
 wire \wave_gen_inst/_0625_ ;
 wire \wave_gen_inst/_0626_ ;
 wire \wave_gen_inst/_0627_ ;
 wire \wave_gen_inst/_0628_ ;
 wire \wave_gen_inst/_0629_ ;
 wire \wave_gen_inst/_0630_ ;
 wire \wave_gen_inst/_0631_ ;
 wire \wave_gen_inst/_0632_ ;
 wire \wave_gen_inst/_0633_ ;
 wire \wave_gen_inst/_0634_ ;
 wire \wave_gen_inst/_0635_ ;
 wire \wave_gen_inst/_0636_ ;
 wire \wave_gen_inst/_0637_ ;
 wire \wave_gen_inst/_0638_ ;
 wire \wave_gen_inst/_0639_ ;
 wire net82;
 wire \wave_gen_inst/_0641_ ;
 wire \wave_gen_inst/_0642_ ;
 wire \wave_gen_inst/_0643_ ;
 wire \wave_gen_inst/_0644_ ;
 wire \wave_gen_inst/_0645_ ;
 wire \wave_gen_inst/_0646_ ;
 wire \wave_gen_inst/_0647_ ;
 wire \wave_gen_inst/_0648_ ;
 wire \wave_gen_inst/_0649_ ;
 wire \wave_gen_inst/_0650_ ;
 wire \wave_gen_inst/_0651_ ;
 wire \wave_gen_inst/_0652_ ;
 wire \wave_gen_inst/_0653_ ;
 wire \wave_gen_inst/_0654_ ;
 wire \wave_gen_inst/_0655_ ;
 wire \wave_gen_inst/_0656_ ;
 wire \wave_gen_inst/_0657_ ;
 wire \wave_gen_inst/_0658_ ;
 wire \wave_gen_inst/_0659_ ;
 wire \wave_gen_inst/_0660_ ;
 wire \wave_gen_inst/_0661_ ;
 wire \wave_gen_inst/_0662_ ;
 wire \wave_gen_inst/_0663_ ;
 wire \wave_gen_inst/_0664_ ;
 wire \wave_gen_inst/_0665_ ;
 wire \wave_gen_inst/_0666_ ;
 wire \wave_gen_inst/_0667_ ;
 wire \wave_gen_inst/_0668_ ;
 wire \wave_gen_inst/_0669_ ;
 wire \wave_gen_inst/_0670_ ;
 wire \wave_gen_inst/_0671_ ;
 wire \wave_gen_inst/_0672_ ;
 wire \wave_gen_inst/_0673_ ;
 wire \wave_gen_inst/_0674_ ;
 wire \wave_gen_inst/_0675_ ;
 wire \wave_gen_inst/_0676_ ;
 wire \wave_gen_inst/_0677_ ;
 wire \wave_gen_inst/_0678_ ;
 wire \wave_gen_inst/_0679_ ;
 wire \wave_gen_inst/_0680_ ;
 wire \wave_gen_inst/_0681_ ;
 wire \wave_gen_inst/_0682_ ;
 wire \wave_gen_inst/_0683_ ;
 wire net81;
 wire \wave_gen_inst/_0685_ ;
 wire \wave_gen_inst/_0686_ ;
 wire \wave_gen_inst/_0687_ ;
 wire \wave_gen_inst/_0688_ ;
 wire \wave_gen_inst/_0689_ ;
 wire \wave_gen_inst/_0690_ ;
 wire \wave_gen_inst/_0691_ ;
 wire \wave_gen_inst/_0692_ ;
 wire \wave_gen_inst/_0693_ ;
 wire \wave_gen_inst/_0694_ ;
 wire \wave_gen_inst/_0695_ ;
 wire \wave_gen_inst/_0696_ ;
 wire \wave_gen_inst/_0697_ ;
 wire \wave_gen_inst/_0698_ ;
 wire \wave_gen_inst/_0699_ ;
 wire \wave_gen_inst/_0700_ ;
 wire \wave_gen_inst/_0701_ ;
 wire \wave_gen_inst/_0702_ ;
 wire \wave_gen_inst/_0703_ ;
 wire \wave_gen_inst/_0704_ ;
 wire \wave_gen_inst/_0705_ ;
 wire \wave_gen_inst/_0706_ ;
 wire \wave_gen_inst/_0707_ ;
 wire \wave_gen_inst/_0708_ ;
 wire \wave_gen_inst/_0709_ ;
 wire \wave_gen_inst/_0710_ ;
 wire \wave_gen_inst/_0711_ ;
 wire \wave_gen_inst/_0712_ ;
 wire \wave_gen_inst/_0713_ ;
 wire \wave_gen_inst/_0714_ ;
 wire \wave_gen_inst/_0715_ ;
 wire \wave_gen_inst/_0716_ ;
 wire \wave_gen_inst/_0717_ ;
 wire \wave_gen_inst/_0718_ ;
 wire net80;
 wire \wave_gen_inst/_0720_ ;
 wire \wave_gen_inst/_0721_ ;
 wire \wave_gen_inst/_0722_ ;
 wire \wave_gen_inst/_0723_ ;
 wire \wave_gen_inst/_0724_ ;
 wire \wave_gen_inst/_0725_ ;
 wire \wave_gen_inst/_0726_ ;
 wire \wave_gen_inst/_0727_ ;
 wire \wave_gen_inst/_0728_ ;
 wire \wave_gen_inst/_0729_ ;
 wire \wave_gen_inst/_0730_ ;
 wire \wave_gen_inst/_0731_ ;
 wire \wave_gen_inst/_0732_ ;
 wire \wave_gen_inst/_0733_ ;
 wire \wave_gen_inst/_0734_ ;
 wire \wave_gen_inst/_0735_ ;
 wire \wave_gen_inst/_0736_ ;
 wire \wave_gen_inst/_0737_ ;
 wire \wave_gen_inst/_0738_ ;
 wire \wave_gen_inst/_0739_ ;
 wire \wave_gen_inst/_0740_ ;
 wire \wave_gen_inst/_0741_ ;
 wire net79;
 wire \wave_gen_inst/_0743_ ;
 wire \wave_gen_inst/_0744_ ;
 wire \wave_gen_inst/_0745_ ;
 wire \wave_gen_inst/_0746_ ;
 wire \wave_gen_inst/_0747_ ;
 wire \wave_gen_inst/_0748_ ;
 wire \wave_gen_inst/_0749_ ;
 wire \wave_gen_inst/_0750_ ;
 wire \wave_gen_inst/_0751_ ;
 wire \wave_gen_inst/_0752_ ;
 wire \wave_gen_inst/_0753_ ;
 wire \wave_gen_inst/_0754_ ;
 wire \wave_gen_inst/_0755_ ;
 wire \wave_gen_inst/_0756_ ;
 wire \wave_gen_inst/_0757_ ;
 wire \wave_gen_inst/_0758_ ;
 wire \wave_gen_inst/_0759_ ;
 wire \wave_gen_inst/_0760_ ;
 wire \wave_gen_inst/_0761_ ;
 wire \wave_gen_inst/_0762_ ;
 wire \wave_gen_inst/_0763_ ;
 wire \wave_gen_inst/_0764_ ;
 wire \wave_gen_inst/_0765_ ;
 wire \wave_gen_inst/_0766_ ;
 wire \wave_gen_inst/_0767_ ;
 wire \wave_gen_inst/_0768_ ;
 wire \wave_gen_inst/_0769_ ;
 wire \wave_gen_inst/_0770_ ;
 wire \wave_gen_inst/_0771_ ;
 wire \wave_gen_inst/_0772_ ;
 wire \wave_gen_inst/_0773_ ;
 wire \wave_gen_inst/_0774_ ;
 wire \wave_gen_inst/_0775_ ;
 wire \wave_gen_inst/_0776_ ;
 wire \wave_gen_inst/_0777_ ;
 wire \wave_gen_inst/_0778_ ;
 wire \wave_gen_inst/_0779_ ;
 wire \wave_gen_inst/_0780_ ;
 wire \wave_gen_inst/_0781_ ;
 wire \wave_gen_inst/_0782_ ;
 wire \wave_gen_inst/_0783_ ;
 wire \wave_gen_inst/_0784_ ;
 wire \wave_gen_inst/_0785_ ;
 wire \wave_gen_inst/_0786_ ;
 wire \wave_gen_inst/_0787_ ;
 wire \wave_gen_inst/_0788_ ;
 wire \wave_gen_inst/_0789_ ;
 wire \wave_gen_inst/_0790_ ;
 wire \wave_gen_inst/_0791_ ;
 wire \wave_gen_inst/_0792_ ;
 wire \wave_gen_inst/_0793_ ;
 wire \wave_gen_inst/_0794_ ;
 wire \wave_gen_inst/_0795_ ;
 wire \wave_gen_inst/_0796_ ;
 wire \wave_gen_inst/_0797_ ;
 wire \wave_gen_inst/_0798_ ;
 wire \wave_gen_inst/_0799_ ;
 wire \wave_gen_inst/_0800_ ;
 wire \wave_gen_inst/_0801_ ;
 wire \wave_gen_inst/_0802_ ;
 wire \wave_gen_inst/_0803_ ;
 wire \wave_gen_inst/_0804_ ;
 wire \wave_gen_inst/_0805_ ;
 wire \wave_gen_inst/_0806_ ;
 wire \wave_gen_inst/_0807_ ;
 wire \wave_gen_inst/_0808_ ;
 wire \wave_gen_inst/_0809_ ;
 wire \wave_gen_inst/_0810_ ;
 wire \wave_gen_inst/_0811_ ;
 wire \wave_gen_inst/_0812_ ;
 wire \wave_gen_inst/_0813_ ;
 wire \wave_gen_inst/_0814_ ;
 wire \wave_gen_inst/_0815_ ;
 wire \wave_gen_inst/_0816_ ;
 wire \wave_gen_inst/_0817_ ;
 wire \wave_gen_inst/_0818_ ;
 wire \wave_gen_inst/_0819_ ;
 wire \wave_gen_inst/_0820_ ;
 wire \wave_gen_inst/_0821_ ;
 wire \wave_gen_inst/_0822_ ;
 wire net78;
 wire net77;
 wire \wave_gen_inst/_0825_ ;
 wire \wave_gen_inst/_0826_ ;
 wire net76;
 wire net75;
 wire \wave_gen_inst/_0829_ ;
 wire net74;
 wire \wave_gen_inst/_0831_ ;
 wire \wave_gen_inst/_0832_ ;
 wire \wave_gen_inst/_0833_ ;
 wire net73;
 wire net72;
 wire \wave_gen_inst/_0836_ ;
 wire \wave_gen_inst/_0837_ ;
 wire \wave_gen_inst/_0838_ ;
 wire \wave_gen_inst/_0839_ ;
 wire \wave_gen_inst/_0840_ ;
 wire \wave_gen_inst/_0841_ ;
 wire \wave_gen_inst/_0842_ ;
 wire \wave_gen_inst/_0843_ ;
 wire \wave_gen_inst/_0844_ ;
 wire \wave_gen_inst/_0845_ ;
 wire \wave_gen_inst/_0846_ ;
 wire \wave_gen_inst/_0847_ ;
 wire \wave_gen_inst/_0848_ ;
 wire \wave_gen_inst/_0849_ ;
 wire \wave_gen_inst/_0850_ ;
 wire \wave_gen_inst/_0851_ ;
 wire \wave_gen_inst/_0852_ ;
 wire \wave_gen_inst/_0853_ ;
 wire \wave_gen_inst/_0854_ ;
 wire \wave_gen_inst/_0855_ ;
 wire \wave_gen_inst/_0856_ ;
 wire \wave_gen_inst/_0857_ ;
 wire \wave_gen_inst/_0858_ ;
 wire \wave_gen_inst/_0859_ ;
 wire \wave_gen_inst/_0860_ ;
 wire \wave_gen_inst/_0861_ ;
 wire \wave_gen_inst/_0862_ ;
 wire \wave_gen_inst/_0863_ ;
 wire \wave_gen_inst/_0864_ ;
 wire \wave_gen_inst/_0865_ ;
 wire \wave_gen_inst/_0866_ ;
 wire \wave_gen_inst/_0867_ ;
 wire \wave_gen_inst/_0868_ ;
 wire \wave_gen_inst/_0869_ ;
 wire \wave_gen_inst/_0870_ ;
 wire \wave_gen_inst/_0871_ ;
 wire \wave_gen_inst/_0872_ ;
 wire \wave_gen_inst/_0873_ ;
 wire \wave_gen_inst/_0874_ ;
 wire \wave_gen_inst/_0875_ ;
 wire \wave_gen_inst/_0876_ ;
 wire \wave_gen_inst/_0877_ ;
 wire \wave_gen_inst/_0878_ ;
 wire \wave_gen_inst/_0879_ ;
 wire \wave_gen_inst/_0880_ ;
 wire \wave_gen_inst/_0881_ ;
 wire \wave_gen_inst/_0882_ ;
 wire \wave_gen_inst/_0883_ ;
 wire \wave_gen_inst/_0884_ ;
 wire \wave_gen_inst/_0885_ ;
 wire \wave_gen_inst/_0886_ ;
 wire \wave_gen_inst/_0887_ ;
 wire \wave_gen_inst/_0888_ ;
 wire \wave_gen_inst/_0889_ ;
 wire \wave_gen_inst/_0890_ ;
 wire \wave_gen_inst/_0891_ ;
 wire \wave_gen_inst/_0892_ ;
 wire \wave_gen_inst/_0893_ ;
 wire \wave_gen_inst/_0894_ ;
 wire \wave_gen_inst/_0895_ ;
 wire \wave_gen_inst/_0896_ ;
 wire \wave_gen_inst/_0897_ ;
 wire \wave_gen_inst/_0898_ ;
 wire \wave_gen_inst/_0899_ ;
 wire \wave_gen_inst/_0900_ ;
 wire \wave_gen_inst/_0901_ ;
 wire \wave_gen_inst/_0902_ ;
 wire \wave_gen_inst/_0903_ ;
 wire \wave_gen_inst/_0904_ ;
 wire \wave_gen_inst/_0905_ ;
 wire \wave_gen_inst/_0906_ ;
 wire \wave_gen_inst/_0907_ ;
 wire \wave_gen_inst/_0908_ ;
 wire \wave_gen_inst/_0909_ ;
 wire \wave_gen_inst/_0910_ ;
 wire \wave_gen_inst/_0911_ ;
 wire \wave_gen_inst/_0912_ ;
 wire \wave_gen_inst/_0913_ ;
 wire \wave_gen_inst/_0914_ ;
 wire \wave_gen_inst/_0915_ ;
 wire \wave_gen_inst/_0916_ ;
 wire \wave_gen_inst/_0917_ ;
 wire \wave_gen_inst/_0918_ ;
 wire \wave_gen_inst/_0919_ ;
 wire \wave_gen_inst/_0920_ ;
 wire \wave_gen_inst/_0921_ ;
 wire net71;
 wire net70;
 wire net69;
 wire \wave_gen_inst/_0925_ ;
 wire \wave_gen_inst/_0926_ ;
 wire \wave_gen_inst/_0927_ ;
 wire net68;
 wire \wave_gen_inst/_0929_ ;
 wire \wave_gen_inst/_0930_ ;
 wire \wave_gen_inst/_0931_ ;
 wire \wave_gen_inst/_0932_ ;
 wire net67;
 wire \wave_gen_inst/_0934_ ;
 wire \wave_gen_inst/_0935_ ;
 wire \wave_gen_inst/_0936_ ;
 wire \wave_gen_inst/_0937_ ;
 wire \wave_gen_inst/_0938_ ;
 wire net66;
 wire \wave_gen_inst/_0940_ ;
 wire \wave_gen_inst/_0941_ ;
 wire \wave_gen_inst/_0942_ ;
 wire \wave_gen_inst/_0943_ ;
 wire \wave_gen_inst/_0944_ ;
 wire \wave_gen_inst/_0945_ ;
 wire \wave_gen_inst/_0946_ ;
 wire \wave_gen_inst/_0947_ ;
 wire \wave_gen_inst/_0948_ ;
 wire net65;
 wire \wave_gen_inst/_0950_ ;
 wire \wave_gen_inst/_0951_ ;
 wire \wave_gen_inst/_0952_ ;
 wire \wave_gen_inst/_0953_ ;
 wire \wave_gen_inst/_0954_ ;
 wire \wave_gen_inst/_0955_ ;
 wire \wave_gen_inst/_0956_ ;
 wire \wave_gen_inst/_0957_ ;
 wire \wave_gen_inst/_0958_ ;
 wire \wave_gen_inst/_0959_ ;
 wire \wave_gen_inst/_0960_ ;
 wire \wave_gen_inst/_0961_ ;
 wire net64;
 wire \wave_gen_inst/_0963_ ;
 wire \wave_gen_inst/_0964_ ;
 wire \wave_gen_inst/_0965_ ;
 wire \wave_gen_inst/_0966_ ;
 wire \wave_gen_inst/_0967_ ;
 wire \wave_gen_inst/_0968_ ;
 wire \wave_gen_inst/_0969_ ;
 wire \wave_gen_inst/_0970_ ;
 wire \wave_gen_inst/_0971_ ;
 wire \wave_gen_inst/_0972_ ;
 wire \wave_gen_inst/_0973_ ;
 wire \wave_gen_inst/_0974_ ;
 wire \wave_gen_inst/_0975_ ;
 wire \wave_gen_inst/_0976_ ;
 wire \wave_gen_inst/_0977_ ;
 wire \wave_gen_inst/_0978_ ;
 wire \wave_gen_inst/_0979_ ;
 wire \wave_gen_inst/_0980_ ;
 wire \wave_gen_inst/_0981_ ;
 wire \wave_gen_inst/_0982_ ;
 wire \wave_gen_inst/_0983_ ;
 wire \wave_gen_inst/_0984_ ;
 wire \wave_gen_inst/_0985_ ;
 wire \wave_gen_inst/_0986_ ;
 wire \wave_gen_inst/_0987_ ;
 wire \wave_gen_inst/_0988_ ;
 wire \wave_gen_inst/_0989_ ;
 wire \wave_gen_inst/_0990_ ;
 wire \wave_gen_inst/_0991_ ;
 wire \wave_gen_inst/_0992_ ;
 wire \wave_gen_inst/_0993_ ;
 wire \wave_gen_inst/_0994_ ;
 wire \wave_gen_inst/_0995_ ;
 wire \wave_gen_inst/_0996_ ;
 wire \wave_gen_inst/_0997_ ;
 wire \wave_gen_inst/_0998_ ;
 wire \wave_gen_inst/_0999_ ;
 wire \wave_gen_inst/_1000_ ;
 wire \wave_gen_inst/_1001_ ;
 wire \wave_gen_inst/_1002_ ;
 wire \wave_gen_inst/_1003_ ;
 wire \wave_gen_inst/_1004_ ;
 wire \wave_gen_inst/_1005_ ;
 wire \wave_gen_inst/_1006_ ;
 wire \wave_gen_inst/_1007_ ;
 wire \wave_gen_inst/_1008_ ;
 wire \wave_gen_inst/_1009_ ;
 wire \wave_gen_inst/_1010_ ;
 wire \wave_gen_inst/_1011_ ;
 wire \wave_gen_inst/_1012_ ;
 wire \wave_gen_inst/_1013_ ;
 wire \wave_gen_inst/_1014_ ;
 wire \wave_gen_inst/_1015_ ;
 wire \wave_gen_inst/_1016_ ;
 wire \wave_gen_inst/_1017_ ;
 wire \wave_gen_inst/_1018_ ;
 wire \wave_gen_inst/_1019_ ;
 wire \wave_gen_inst/_1020_ ;
 wire \wave_gen_inst/_1021_ ;
 wire \wave_gen_inst/_1022_ ;
 wire \wave_gen_inst/_1023_ ;
 wire \wave_gen_inst/_1024_ ;
 wire \wave_gen_inst/_1025_ ;
 wire \wave_gen_inst/_1026_ ;
 wire \wave_gen_inst/_1027_ ;
 wire \wave_gen_inst/_1028_ ;
 wire \wave_gen_inst/_1029_ ;
 wire \wave_gen_inst/_1030_ ;
 wire \wave_gen_inst/_1031_ ;
 wire net63;
 wire \wave_gen_inst/_1033_ ;
 wire \wave_gen_inst/_1034_ ;
 wire \wave_gen_inst/_1035_ ;
 wire \wave_gen_inst/_1036_ ;
 wire \wave_gen_inst/_1037_ ;
 wire \wave_gen_inst/_1038_ ;
 wire \wave_gen_inst/_1039_ ;
 wire \wave_gen_inst/_1040_ ;
 wire \wave_gen_inst/_1041_ ;
 wire \wave_gen_inst/_1042_ ;
 wire \wave_gen_inst/_1043_ ;
 wire \wave_gen_inst/_1044_ ;
 wire \wave_gen_inst/_1045_ ;
 wire \wave_gen_inst/_1046_ ;
 wire \wave_gen_inst/_1047_ ;
 wire \wave_gen_inst/_1048_ ;
 wire \wave_gen_inst/_1049_ ;
 wire \wave_gen_inst/_1050_ ;
 wire \wave_gen_inst/_1051_ ;
 wire \wave_gen_inst/_1052_ ;
 wire \wave_gen_inst/_1053_ ;
 wire \wave_gen_inst/_1054_ ;
 wire \wave_gen_inst/_1055_ ;
 wire \wave_gen_inst/_1056_ ;
 wire \wave_gen_inst/_1057_ ;
 wire \wave_gen_inst/_1058_ ;
 wire \wave_gen_inst/_1059_ ;
 wire \wave_gen_inst/_1060_ ;
 wire \wave_gen_inst/_1061_ ;
 wire \wave_gen_inst/_1062_ ;
 wire \wave_gen_inst/_1063_ ;
 wire \wave_gen_inst/_1064_ ;
 wire \wave_gen_inst/_1065_ ;
 wire net62;
 wire \wave_gen_inst/_1067_ ;
 wire \wave_gen_inst/_1068_ ;
 wire \wave_gen_inst/_1069_ ;
 wire \wave_gen_inst/_1070_ ;
 wire \wave_gen_inst/_1071_ ;
 wire \wave_gen_inst/_1072_ ;
 wire \wave_gen_inst/_1073_ ;
 wire \wave_gen_inst/_1074_ ;
 wire \wave_gen_inst/_1075_ ;
 wire \wave_gen_inst/_1076_ ;
 wire \wave_gen_inst/_1077_ ;
 wire \wave_gen_inst/_1078_ ;
 wire \wave_gen_inst/_1079_ ;
 wire \wave_gen_inst/_1080_ ;
 wire \wave_gen_inst/_1081_ ;
 wire \wave_gen_inst/_1082_ ;
 wire \wave_gen_inst/_1083_ ;
 wire \wave_gen_inst/_1084_ ;
 wire \wave_gen_inst/_1085_ ;
 wire \wave_gen_inst/_1086_ ;
 wire \wave_gen_inst/_1087_ ;
 wire \wave_gen_inst/_1088_ ;
 wire \wave_gen_inst/_1089_ ;
 wire \wave_gen_inst/_1090_ ;
 wire \wave_gen_inst/_1091_ ;
 wire \wave_gen_inst/_1092_ ;
 wire net61;
 wire \wave_gen_inst/_1094_ ;
 wire \wave_gen_inst/_1095_ ;
 wire \wave_gen_inst/_1096_ ;
 wire \wave_gen_inst/_1097_ ;
 wire \wave_gen_inst/_1098_ ;
 wire \wave_gen_inst/_1099_ ;
 wire net60;
 wire \wave_gen_inst/_1101_ ;
 wire \wave_gen_inst/_1102_ ;
 wire \wave_gen_inst/_1103_ ;
 wire \wave_gen_inst/_1104_ ;
 wire \wave_gen_inst/_1105_ ;
 wire \wave_gen_inst/_1106_ ;
 wire \wave_gen_inst/_1107_ ;
 wire \wave_gen_inst/_1108_ ;
 wire \wave_gen_inst/_1109_ ;
 wire \wave_gen_inst/_1110_ ;
 wire \wave_gen_inst/_1111_ ;
 wire \wave_gen_inst/_1112_ ;
 wire \wave_gen_inst/_1113_ ;
 wire \wave_gen_inst/_1114_ ;
 wire \wave_gen_inst/_1115_ ;
 wire \wave_gen_inst/_1116_ ;
 wire \wave_gen_inst/_1117_ ;
 wire \wave_gen_inst/_1118_ ;
 wire \wave_gen_inst/_1119_ ;
 wire \wave_gen_inst/_1120_ ;
 wire net59;
 wire \wave_gen_inst/_1122_ ;
 wire \wave_gen_inst/_1123_ ;
 wire \wave_gen_inst/_1124_ ;
 wire \wave_gen_inst/_1125_ ;
 wire \wave_gen_inst/_1126_ ;
 wire \wave_gen_inst/_1127_ ;
 wire \wave_gen_inst/_1128_ ;
 wire \wave_gen_inst/_1129_ ;
 wire \wave_gen_inst/_1130_ ;
 wire \wave_gen_inst/_1131_ ;
 wire \wave_gen_inst/_1132_ ;
 wire \wave_gen_inst/_1133_ ;
 wire \wave_gen_inst/_1134_ ;
 wire \wave_gen_inst/_1135_ ;
 wire \wave_gen_inst/_1136_ ;
 wire \wave_gen_inst/_1137_ ;
 wire \wave_gen_inst/_1138_ ;
 wire \wave_gen_inst/_1139_ ;
 wire \wave_gen_inst/_1140_ ;
 wire \wave_gen_inst/_1141_ ;
 wire \wave_gen_inst/_1142_ ;
 wire \wave_gen_inst/_1143_ ;
 wire \wave_gen_inst/_1144_ ;
 wire \wave_gen_inst/_1145_ ;
 wire \wave_gen_inst/_1146_ ;
 wire \wave_gen_inst/_1147_ ;
 wire \wave_gen_inst/_1148_ ;
 wire \wave_gen_inst/_1149_ ;
 wire \wave_gen_inst/_1150_ ;
 wire \wave_gen_inst/_1151_ ;
 wire \wave_gen_inst/_1152_ ;
 wire \wave_gen_inst/_1153_ ;
 wire \wave_gen_inst/_1154_ ;
 wire \wave_gen_inst/_1155_ ;
 wire \wave_gen_inst/_1156_ ;
 wire \wave_gen_inst/_1157_ ;
 wire \wave_gen_inst/_1158_ ;
 wire \wave_gen_inst/_1159_ ;
 wire \wave_gen_inst/_1160_ ;
 wire \wave_gen_inst/_1161_ ;
 wire \wave_gen_inst/_1162_ ;
 wire \wave_gen_inst/_1163_ ;
 wire \wave_gen_inst/_1164_ ;
 wire \wave_gen_inst/_1165_ ;
 wire \wave_gen_inst/_1166_ ;
 wire \wave_gen_inst/_1167_ ;
 wire \wave_gen_inst/_1168_ ;
 wire \wave_gen_inst/_1169_ ;
 wire \wave_gen_inst/_1170_ ;
 wire \wave_gen_inst/_1171_ ;
 wire net58;
 wire \wave_gen_inst/_1173_ ;
 wire \wave_gen_inst/_1174_ ;
 wire \wave_gen_inst/_1175_ ;
 wire \wave_gen_inst/_1176_ ;
 wire \wave_gen_inst/_1177_ ;
 wire \wave_gen_inst/_1178_ ;
 wire \wave_gen_inst/_1179_ ;
 wire \wave_gen_inst/_1180_ ;
 wire \wave_gen_inst/_1181_ ;
 wire \wave_gen_inst/_1182_ ;
 wire \wave_gen_inst/_1183_ ;
 wire \wave_gen_inst/_1184_ ;
 wire \wave_gen_inst/_1185_ ;
 wire \wave_gen_inst/_1186_ ;
 wire \wave_gen_inst/_1187_ ;
 wire \wave_gen_inst/_1188_ ;
 wire \wave_gen_inst/_1189_ ;
 wire \wave_gen_inst/_1190_ ;
 wire \wave_gen_inst/_1191_ ;
 wire \wave_gen_inst/_1192_ ;
 wire \wave_gen_inst/_1193_ ;
 wire \wave_gen_inst/_1194_ ;
 wire \wave_gen_inst/_1195_ ;
 wire \wave_gen_inst/_1196_ ;
 wire \wave_gen_inst/_1197_ ;
 wire \wave_gen_inst/_1198_ ;
 wire \wave_gen_inst/_1199_ ;
 wire \wave_gen_inst/_1200_ ;
 wire \wave_gen_inst/_1201_ ;
 wire \wave_gen_inst/_1202_ ;
 wire \wave_gen_inst/_1203_ ;
 wire \wave_gen_inst/_1204_ ;
 wire \wave_gen_inst/_1205_ ;
 wire \wave_gen_inst/_1206_ ;
 wire \wave_gen_inst/_1207_ ;
 wire \wave_gen_inst/_1208_ ;
 wire \wave_gen_inst/_1209_ ;
 wire \wave_gen_inst/_1210_ ;
 wire \wave_gen_inst/_1211_ ;
 wire \wave_gen_inst/_1212_ ;
 wire \wave_gen_inst/_1213_ ;
 wire \wave_gen_inst/_1214_ ;
 wire \wave_gen_inst/_1215_ ;
 wire \wave_gen_inst/_1216_ ;
 wire \wave_gen_inst/_1217_ ;
 wire \wave_gen_inst/_1218_ ;
 wire \wave_gen_inst/_1219_ ;
 wire \wave_gen_inst/_1220_ ;
 wire \wave_gen_inst/_1221_ ;
 wire \wave_gen_inst/_1222_ ;
 wire \wave_gen_inst/_1223_ ;
 wire \wave_gen_inst/_1224_ ;
 wire \wave_gen_inst/_1225_ ;
 wire \wave_gen_inst/_1226_ ;
 wire \wave_gen_inst/_1227_ ;
 wire \wave_gen_inst/_1228_ ;
 wire \wave_gen_inst/_1229_ ;
 wire \wave_gen_inst/_1230_ ;
 wire \wave_gen_inst/_1231_ ;
 wire \wave_gen_inst/_1232_ ;
 wire \wave_gen_inst/_1233_ ;
 wire \wave_gen_inst/_1234_ ;
 wire \wave_gen_inst/_1235_ ;
 wire \wave_gen_inst/_1236_ ;
 wire \wave_gen_inst/_1237_ ;
 wire \wave_gen_inst/_1238_ ;
 wire \wave_gen_inst/_1239_ ;
 wire \wave_gen_inst/_1240_ ;
 wire \wave_gen_inst/_1241_ ;
 wire \wave_gen_inst/_1242_ ;
 wire \wave_gen_inst/_1243_ ;
 wire \wave_gen_inst/_1244_ ;
 wire \wave_gen_inst/_1245_ ;
 wire \wave_gen_inst/_1246_ ;
 wire \wave_gen_inst/_1247_ ;
 wire \wave_gen_inst/_1248_ ;
 wire \wave_gen_inst/_1249_ ;
 wire \wave_gen_inst/_1250_ ;
 wire \wave_gen_inst/_1251_ ;
 wire \wave_gen_inst/_1252_ ;
 wire \wave_gen_inst/_1253_ ;
 wire \wave_gen_inst/_1254_ ;
 wire \wave_gen_inst/_1255_ ;
 wire \wave_gen_inst/_1256_ ;
 wire \wave_gen_inst/_1257_ ;
 wire \wave_gen_inst/_1258_ ;
 wire \wave_gen_inst/_1259_ ;
 wire \wave_gen_inst/_1260_ ;
 wire \wave_gen_inst/_1261_ ;
 wire \wave_gen_inst/_1262_ ;
 wire \wave_gen_inst/_1263_ ;
 wire \wave_gen_inst/_1264_ ;
 wire \wave_gen_inst/_1265_ ;
 wire \wave_gen_inst/_1266_ ;
 wire \wave_gen_inst/_1267_ ;
 wire \wave_gen_inst/_1268_ ;
 wire \wave_gen_inst/_1269_ ;
 wire \wave_gen_inst/_1270_ ;
 wire \wave_gen_inst/_1271_ ;
 wire \wave_gen_inst/_1272_ ;
 wire \wave_gen_inst/_1273_ ;
 wire \wave_gen_inst/_1274_ ;
 wire \wave_gen_inst/_1275_ ;
 wire \wave_gen_inst/_1276_ ;
 wire \wave_gen_inst/_1277_ ;
 wire \wave_gen_inst/_1278_ ;
 wire \wave_gen_inst/_1279_ ;
 wire \wave_gen_inst/_1280_ ;
 wire \wave_gen_inst/_1281_ ;
 wire \wave_gen_inst/_1282_ ;
 wire \wave_gen_inst/_1283_ ;
 wire \wave_gen_inst/_1284_ ;
 wire \wave_gen_inst/_1285_ ;
 wire \wave_gen_inst/_1286_ ;
 wire \wave_gen_inst/_1287_ ;
 wire \wave_gen_inst/_1288_ ;
 wire \wave_gen_inst/_1289_ ;
 wire \wave_gen_inst/_1290_ ;
 wire \wave_gen_inst/_1291_ ;
 wire \wave_gen_inst/_1292_ ;
 wire \wave_gen_inst/_1293_ ;
 wire \wave_gen_inst/_1294_ ;
 wire \wave_gen_inst/_1295_ ;
 wire \wave_gen_inst/_1296_ ;
 wire \wave_gen_inst/_1297_ ;
 wire \wave_gen_inst/_1298_ ;
 wire \wave_gen_inst/_1299_ ;
 wire \wave_gen_inst/_1300_ ;
 wire \wave_gen_inst/_1301_ ;
 wire \wave_gen_inst/_1302_ ;
 wire \wave_gen_inst/_1303_ ;
 wire \wave_gen_inst/_1304_ ;
 wire \wave_gen_inst/_1305_ ;
 wire \wave_gen_inst/_1306_ ;
 wire \wave_gen_inst/_1307_ ;
 wire \wave_gen_inst/_1308_ ;
 wire \wave_gen_inst/_1309_ ;
 wire \wave_gen_inst/_1310_ ;
 wire \wave_gen_inst/_1311_ ;
 wire \wave_gen_inst/_1312_ ;
 wire \wave_gen_inst/_1313_ ;
 wire \wave_gen_inst/_1314_ ;
 wire \wave_gen_inst/_1315_ ;
 wire \wave_gen_inst/_1316_ ;
 wire \wave_gen_inst/_1317_ ;
 wire \wave_gen_inst/_1318_ ;
 wire \wave_gen_inst/_1319_ ;
 wire \wave_gen_inst/_1320_ ;
 wire \wave_gen_inst/_1321_ ;
 wire \wave_gen_inst/_1322_ ;
 wire \wave_gen_inst/_1323_ ;
 wire \wave_gen_inst/_1324_ ;
 wire \wave_gen_inst/_1325_ ;
 wire \wave_gen_inst/_1326_ ;
 wire \wave_gen_inst/_1327_ ;
 wire \wave_gen_inst/_1328_ ;
 wire \wave_gen_inst/_1329_ ;
 wire \wave_gen_inst/_1330_ ;
 wire \wave_gen_inst/_1331_ ;
 wire \wave_gen_inst/_1332_ ;
 wire \wave_gen_inst/_1333_ ;
 wire \wave_gen_inst/_1334_ ;
 wire \wave_gen_inst/_1335_ ;
 wire \wave_gen_inst/_1336_ ;
 wire \wave_gen_inst/_1337_ ;
 wire \wave_gen_inst/_1338_ ;
 wire \wave_gen_inst/_1339_ ;
 wire \wave_gen_inst/_1340_ ;
 wire \wave_gen_inst/_1341_ ;
 wire \wave_gen_inst/_1342_ ;
 wire \wave_gen_inst/_1343_ ;
 wire \wave_gen_inst/_1344_ ;
 wire \wave_gen_inst/_1345_ ;
 wire \wave_gen_inst/_1346_ ;
 wire \wave_gen_inst/_1347_ ;
 wire \wave_gen_inst/_1348_ ;
 wire \wave_gen_inst/_1349_ ;
 wire \wave_gen_inst/_1350_ ;
 wire \wave_gen_inst/_1351_ ;
 wire \wave_gen_inst/_1352_ ;
 wire \wave_gen_inst/_1353_ ;
 wire \wave_gen_inst/_1354_ ;
 wire \wave_gen_inst/_1355_ ;
 wire \wave_gen_inst/_1356_ ;
 wire \wave_gen_inst/_1357_ ;
 wire \wave_gen_inst/_1358_ ;
 wire \wave_gen_inst/_1359_ ;
 wire \wave_gen_inst/_1360_ ;
 wire \wave_gen_inst/_1361_ ;
 wire \wave_gen_inst/_1362_ ;
 wire \wave_gen_inst/_1363_ ;
 wire \wave_gen_inst/_1364_ ;
 wire \wave_gen_inst/_1365_ ;
 wire \wave_gen_inst/_1366_ ;
 wire \wave_gen_inst/_1367_ ;
 wire \wave_gen_inst/_1368_ ;
 wire \wave_gen_inst/_1369_ ;
 wire \wave_gen_inst/_1370_ ;
 wire \wave_gen_inst/_1371_ ;
 wire \wave_gen_inst/_1372_ ;
 wire \wave_gen_inst/_1373_ ;
 wire \wave_gen_inst/_1374_ ;
 wire \wave_gen_inst/_1375_ ;
 wire \wave_gen_inst/_1376_ ;
 wire \wave_gen_inst/_1377_ ;
 wire \wave_gen_inst/_1378_ ;
 wire \wave_gen_inst/_1379_ ;
 wire \wave_gen_inst/_1380_ ;
 wire \wave_gen_inst/_1381_ ;
 wire \wave_gen_inst/_1382_ ;
 wire \wave_gen_inst/_1383_ ;
 wire \wave_gen_inst/_1384_ ;
 wire \wave_gen_inst/_1385_ ;
 wire \wave_gen_inst/_1386_ ;
 wire \wave_gen_inst/_1387_ ;
 wire \wave_gen_inst/_1388_ ;
 wire \wave_gen_inst/_1389_ ;
 wire \wave_gen_inst/_1390_ ;
 wire \wave_gen_inst/_1391_ ;
 wire \wave_gen_inst/_1392_ ;
 wire \wave_gen_inst/_1393_ ;
 wire \wave_gen_inst/_1394_ ;
 wire \wave_gen_inst/_1395_ ;
 wire \wave_gen_inst/_1396_ ;
 wire \wave_gen_inst/_1397_ ;
 wire \wave_gen_inst/_1398_ ;
 wire \wave_gen_inst/_1399_ ;
 wire \wave_gen_inst/_1400_ ;
 wire \wave_gen_inst/_1401_ ;
 wire \wave_gen_inst/_1402_ ;
 wire \wave_gen_inst/_1403_ ;
 wire \wave_gen_inst/_1404_ ;
 wire \wave_gen_inst/_1405_ ;
 wire \wave_gen_inst/_1406_ ;
 wire \wave_gen_inst/_1407_ ;
 wire \wave_gen_inst/_1408_ ;
 wire \wave_gen_inst/_1409_ ;
 wire \wave_gen_inst/_1410_ ;
 wire \wave_gen_inst/_1411_ ;
 wire \wave_gen_inst/_1412_ ;
 wire \wave_gen_inst/_1413_ ;
 wire \wave_gen_inst/_1414_ ;
 wire \wave_gen_inst/_1415_ ;
 wire \wave_gen_inst/_1416_ ;
 wire \wave_gen_inst/_1417_ ;
 wire \wave_gen_inst/_1418_ ;
 wire \wave_gen_inst/_1419_ ;
 wire \wave_gen_inst/_1420_ ;
 wire \wave_gen_inst/_1421_ ;
 wire \wave_gen_inst/_1422_ ;
 wire \wave_gen_inst/_1423_ ;
 wire \wave_gen_inst/_1424_ ;
 wire \wave_gen_inst/_1425_ ;
 wire \wave_gen_inst/_1426_ ;
 wire \wave_gen_inst/_1427_ ;
 wire \wave_gen_inst/_1428_ ;
 wire \wave_gen_inst/_1429_ ;
 wire \wave_gen_inst/_1430_ ;
 wire \wave_gen_inst/_1431_ ;
 wire \wave_gen_inst/_1432_ ;
 wire \wave_gen_inst/_1433_ ;
 wire \wave_gen_inst/_1434_ ;
 wire \wave_gen_inst/_1435_ ;
 wire \wave_gen_inst/_1436_ ;
 wire \wave_gen_inst/_1437_ ;
 wire \wave_gen_inst/_1438_ ;
 wire \wave_gen_inst/_1439_ ;
 wire \wave_gen_inst/_1440_ ;
 wire \wave_gen_inst/_1441_ ;
 wire \wave_gen_inst/_1442_ ;
 wire \wave_gen_inst/_1443_ ;
 wire \wave_gen_inst/_1444_ ;
 wire \wave_gen_inst/_1445_ ;
 wire \wave_gen_inst/_1446_ ;
 wire \wave_gen_inst/_1447_ ;
 wire \wave_gen_inst/_1448_ ;
 wire \wave_gen_inst/_1449_ ;
 wire \wave_gen_inst/_1450_ ;
 wire \wave_gen_inst/_1451_ ;
 wire \wave_gen_inst/_1452_ ;
 wire \wave_gen_inst/_1453_ ;
 wire \wave_gen_inst/_1454_ ;
 wire \wave_gen_inst/_1455_ ;
 wire \wave_gen_inst/_1456_ ;
 wire \wave_gen_inst/_1457_ ;
 wire \wave_gen_inst/_1458_ ;
 wire \wave_gen_inst/_1459_ ;
 wire \wave_gen_inst/_1460_ ;
 wire \wave_gen_inst/_1461_ ;
 wire \wave_gen_inst/_1462_ ;
 wire \wave_gen_inst/_1463_ ;
 wire \wave_gen_inst/_1464_ ;
 wire \wave_gen_inst/_1465_ ;
 wire \wave_gen_inst/_1466_ ;
 wire \wave_gen_inst/_1467_ ;
 wire \wave_gen_inst/_1468_ ;
 wire \wave_gen_inst/_1469_ ;
 wire \wave_gen_inst/_1470_ ;
 wire \wave_gen_inst/_1471_ ;
 wire \wave_gen_inst/_1472_ ;
 wire \wave_gen_inst/_1473_ ;
 wire \wave_gen_inst/_1474_ ;
 wire \wave_gen_inst/_1475_ ;
 wire \wave_gen_inst/_1476_ ;
 wire \wave_gen_inst/_1477_ ;
 wire \wave_gen_inst/_1478_ ;
 wire \wave_gen_inst/_1479_ ;
 wire \wave_gen_inst/_1480_ ;
 wire \wave_gen_inst/_1481_ ;
 wire \wave_gen_inst/_1482_ ;
 wire \wave_gen_inst/_1483_ ;
 wire \wave_gen_inst/_1484_ ;
 wire \wave_gen_inst/_1485_ ;
 wire \wave_gen_inst/_1486_ ;
 wire \wave_gen_inst/_1487_ ;
 wire \wave_gen_inst/_1488_ ;
 wire \wave_gen_inst/_1489_ ;
 wire \wave_gen_inst/_1490_ ;
 wire \wave_gen_inst/_1491_ ;
 wire \wave_gen_inst/_1492_ ;
 wire \wave_gen_inst/_1493_ ;
 wire \wave_gen_inst/_1494_ ;
 wire \wave_gen_inst/_1495_ ;
 wire \wave_gen_inst/_1496_ ;
 wire \wave_gen_inst/_1497_ ;
 wire \wave_gen_inst/_1498_ ;
 wire \wave_gen_inst/_1499_ ;
 wire \wave_gen_inst/_1500_ ;
 wire \wave_gen_inst/_1501_ ;
 wire \wave_gen_inst/_1502_ ;
 wire \wave_gen_inst/_1503_ ;
 wire \wave_gen_inst/_1504_ ;
 wire \wave_gen_inst/_1505_ ;
 wire \wave_gen_inst/_1506_ ;
 wire \wave_gen_inst/_1507_ ;
 wire \wave_gen_inst/_1508_ ;
 wire net229;
 wire net228;
 wire net227;
 wire net226;
 wire net225;
 wire \wave_gen_inst/_1514_ ;
 wire net224;
 wire net223;
 wire net222;
 wire net221;
 wire net220;
 wire net219;
 wire net218;
 wire net217;
 wire net216;
 wire net215;
 wire \wave_gen_inst/_1525_ ;
 wire \wave_gen_inst/_1526_ ;
 wire net214;
 wire \wave_gen_inst/_1528_ ;
 wire net213;
 wire net212;
 wire \wave_gen_inst/_1531_ ;
 wire net211;
 wire \wave_gen_inst/_1533_ ;
 wire net210;
 wire \wave_gen_inst/_1535_ ;
 wire net209;
 wire \wave_gen_inst/_1537_ ;
 wire \wave_gen_inst/_1538_ ;
 wire net208;
 wire net207;
 wire \wave_gen_inst/_1541_ ;
 wire net206;
 wire net205;
 wire \wave_gen_inst/_1544_ ;
 wire \wave_gen_inst/_1545_ ;
 wire \wave_gen_inst/_1546_ ;
 wire \wave_gen_inst/_1547_ ;
 wire \wave_gen_inst/_1548_ ;
 wire net204;
 wire \wave_gen_inst/_1550_ ;
 wire \wave_gen_inst/_1551_ ;
 wire \wave_gen_inst/_1552_ ;
 wire net203;
 wire \wave_gen_inst/_1554_ ;
 wire \wave_gen_inst/_1555_ ;
 wire \wave_gen_inst/_1556_ ;
 wire net202;
 wire \wave_gen_inst/_1558_ ;
 wire net201;
 wire net200;
 wire \wave_gen_inst/_1561_ ;
 wire \wave_gen_inst/_1562_ ;
 wire net199;
 wire net198;
 wire net197;
 wire \wave_gen_inst/_1566_ ;
 wire \wave_gen_inst/_1567_ ;
 wire \wave_gen_inst/_1568_ ;
 wire \wave_gen_inst/_1569_ ;
 wire \wave_gen_inst/_1570_ ;
 wire \wave_gen_inst/_1571_ ;
 wire \wave_gen_inst/_1572_ ;
 wire net196;
 wire \wave_gen_inst/_1574_ ;
 wire \wave_gen_inst/_1575_ ;
 wire net195;
 wire net194;
 wire \wave_gen_inst/_1578_ ;
 wire net193;
 wire \wave_gen_inst/_1580_ ;
 wire \wave_gen_inst/_1581_ ;
 wire \wave_gen_inst/_1582_ ;
 wire net192;
 wire net191;
 wire net190;
 wire \wave_gen_inst/_1586_ ;
 wire \wave_gen_inst/_1587_ ;
 wire \wave_gen_inst/_1588_ ;
 wire net189;
 wire \wave_gen_inst/_1590_ ;
 wire net188;
 wire \wave_gen_inst/_1592_ ;
 wire \wave_gen_inst/_1593_ ;
 wire net187;
 wire net186;
 wire \wave_gen_inst/_1596_ ;
 wire \wave_gen_inst/_1597_ ;
 wire \wave_gen_inst/_1598_ ;
 wire \wave_gen_inst/_1599_ ;
 wire \wave_gen_inst/_1600_ ;
 wire \wave_gen_inst/_1601_ ;
 wire \wave_gen_inst/_1602_ ;
 wire net185;
 wire net184;
 wire net183;
 wire \wave_gen_inst/_1606_ ;
 wire \wave_gen_inst/_1607_ ;
 wire \wave_gen_inst/_1608_ ;
 wire net182;
 wire net181;
 wire \wave_gen_inst/_1611_ ;
 wire net180;
 wire \wave_gen_inst/_1613_ ;
 wire \wave_gen_inst/_1614_ ;
 wire \wave_gen_inst/_1615_ ;
 wire \wave_gen_inst/_1616_ ;
 wire net179;
 wire net178;
 wire net177;
 wire \wave_gen_inst/_1620_ ;
 wire net176;
 wire \wave_gen_inst/_1622_ ;
 wire \wave_gen_inst/_1623_ ;
 wire net175;
 wire net174;
 wire net173;
 wire \wave_gen_inst/_1627_ ;
 wire \wave_gen_inst/_1628_ ;
 wire \wave_gen_inst/_1629_ ;
 wire \wave_gen_inst/_1630_ ;
 wire \wave_gen_inst/_1631_ ;
 wire \wave_gen_inst/_1632_ ;
 wire net172;
 wire net171;
 wire \wave_gen_inst/_1635_ ;
 wire \wave_gen_inst/_1636_ ;
 wire \wave_gen_inst/_1637_ ;
 wire \wave_gen_inst/_1638_ ;
 wire \wave_gen_inst/_1639_ ;
 wire \wave_gen_inst/_1640_ ;
 wire \wave_gen_inst/_1641_ ;
 wire \wave_gen_inst/_1642_ ;
 wire \wave_gen_inst/_1643_ ;
 wire \wave_gen_inst/_1644_ ;
 wire \wave_gen_inst/_1645_ ;
 wire \wave_gen_inst/_1646_ ;
 wire net170;
 wire \wave_gen_inst/_1648_ ;
 wire \wave_gen_inst/_1649_ ;
 wire \wave_gen_inst/_1650_ ;
 wire \wave_gen_inst/_1651_ ;
 wire \wave_gen_inst/_1652_ ;
 wire \wave_gen_inst/_1653_ ;
 wire \wave_gen_inst/_1654_ ;
 wire \wave_gen_inst/_1655_ ;
 wire \wave_gen_inst/_1656_ ;
 wire \wave_gen_inst/_1657_ ;
 wire \wave_gen_inst/_1658_ ;
 wire \wave_gen_inst/_1659_ ;
 wire \wave_gen_inst/_1660_ ;
 wire \wave_gen_inst/_1661_ ;
 wire \wave_gen_inst/_1662_ ;
 wire \wave_gen_inst/_1663_ ;
 wire net169;
 wire \wave_gen_inst/_1665_ ;
 wire \wave_gen_inst/_1666_ ;
 wire \wave_gen_inst/_1667_ ;
 wire \wave_gen_inst/_1668_ ;
 wire \wave_gen_inst/_1669_ ;
 wire \wave_gen_inst/_1670_ ;
 wire \wave_gen_inst/_1671_ ;
 wire \wave_gen_inst/_1672_ ;
 wire \wave_gen_inst/_1673_ ;
 wire \wave_gen_inst/_1674_ ;
 wire \wave_gen_inst/_1675_ ;
 wire \wave_gen_inst/_1676_ ;
 wire \wave_gen_inst/_1677_ ;
 wire \wave_gen_inst/_1678_ ;
 wire \wave_gen_inst/_1679_ ;
 wire \wave_gen_inst/_1680_ ;
 wire \wave_gen_inst/_1681_ ;
 wire \wave_gen_inst/_1682_ ;
 wire \wave_gen_inst/_1683_ ;
 wire \wave_gen_inst/_1684_ ;
 wire \wave_gen_inst/_1685_ ;
 wire \wave_gen_inst/_1686_ ;
 wire \wave_gen_inst/_1687_ ;
 wire \wave_gen_inst/_1688_ ;
 wire \wave_gen_inst/_1689_ ;
 wire \wave_gen_inst/_1690_ ;
 wire \wave_gen_inst/_1691_ ;
 wire \wave_gen_inst/_1692_ ;
 wire \wave_gen_inst/_1693_ ;
 wire \wave_gen_inst/_1694_ ;
 wire \wave_gen_inst/_1695_ ;
 wire \wave_gen_inst/_1696_ ;
 wire \wave_gen_inst/_1697_ ;
 wire \wave_gen_inst/_1698_ ;
 wire \wave_gen_inst/_1699_ ;
 wire \wave_gen_inst/_1700_ ;
 wire \wave_gen_inst/_1701_ ;
 wire \wave_gen_inst/_1702_ ;
 wire \wave_gen_inst/_1703_ ;
 wire \wave_gen_inst/_1704_ ;
 wire \wave_gen_inst/_1705_ ;
 wire \wave_gen_inst/_1706_ ;
 wire \wave_gen_inst/_1707_ ;
 wire \wave_gen_inst/_1708_ ;
 wire \wave_gen_inst/_1709_ ;
 wire \wave_gen_inst/_1710_ ;
 wire \wave_gen_inst/_1711_ ;
 wire \wave_gen_inst/_1712_ ;
 wire \wave_gen_inst/_1713_ ;
 wire \wave_gen_inst/_1714_ ;
 wire \wave_gen_inst/_1715_ ;
 wire \wave_gen_inst/_1716_ ;
 wire \wave_gen_inst/_1717_ ;
 wire \wave_gen_inst/_1718_ ;
 wire \wave_gen_inst/_1719_ ;
 wire \wave_gen_inst/_1720_ ;
 wire \wave_gen_inst/_1721_ ;
 wire \wave_gen_inst/_1722_ ;
 wire \wave_gen_inst/_1723_ ;
 wire \wave_gen_inst/_1724_ ;
 wire \wave_gen_inst/_1725_ ;
 wire \wave_gen_inst/_1726_ ;
 wire \wave_gen_inst/_1727_ ;
 wire \wave_gen_inst/_1728_ ;
 wire \wave_gen_inst/_1729_ ;
 wire \wave_gen_inst/_1730_ ;
 wire \wave_gen_inst/_1731_ ;
 wire \wave_gen_inst/_1732_ ;
 wire \wave_gen_inst/_1733_ ;
 wire \wave_gen_inst/_1734_ ;
 wire \wave_gen_inst/_1735_ ;
 wire \wave_gen_inst/_1736_ ;
 wire \wave_gen_inst/_1737_ ;
 wire \wave_gen_inst/_1738_ ;
 wire \wave_gen_inst/_1739_ ;
 wire \wave_gen_inst/_1740_ ;
 wire \wave_gen_inst/_1741_ ;
 wire \wave_gen_inst/_1742_ ;
 wire \wave_gen_inst/_1743_ ;
 wire \wave_gen_inst/_1744_ ;
 wire \wave_gen_inst/_1745_ ;
 wire \wave_gen_inst/_1746_ ;
 wire \wave_gen_inst/_1747_ ;
 wire \wave_gen_inst/_1748_ ;
 wire net168;
 wire net167;
 wire net166;
 wire \wave_gen_inst/_1752_ ;
 wire \wave_gen_inst/_1753_ ;
 wire net165;
 wire \wave_gen_inst/_1755_ ;
 wire net164;
 wire net163;
 wire \wave_gen_inst/_1758_ ;
 wire net162;
 wire net161;
 wire net160;
 wire \wave_gen_inst/_1762_ ;
 wire \wave_gen_inst/_1763_ ;
 wire net159;
 wire net158;
 wire net157;
 wire \wave_gen_inst/_1767_ ;
 wire net156;
 wire net155;
 wire \wave_gen_inst/_1770_ ;
 wire \wave_gen_inst/_1771_ ;
 wire net154;
 wire net153;
 wire \wave_gen_inst/_1774_ ;
 wire net152;
 wire net151;
 wire net150;
 wire \wave_gen_inst/_1778_ ;
 wire \wave_gen_inst/_1779_ ;
 wire \wave_gen_inst/_1780_ ;
 wire net149;
 wire net148;
 wire \wave_gen_inst/_1783_ ;
 wire net147;
 wire net146;
 wire \wave_gen_inst/_1786_ ;
 wire \wave_gen_inst/_1787_ ;
 wire net145;
 wire net144;
 wire \wave_gen_inst/_1790_ ;
 wire net143;
 wire net142;
 wire \wave_gen_inst/_1793_ ;
 wire \wave_gen_inst/_1794_ ;
 wire \wave_gen_inst/_1795_ ;
 wire net141;
 wire net140;
 wire \wave_gen_inst/_1798_ ;
 wire net139;
 wire net138;
 wire \wave_gen_inst/_1801_ ;
 wire \wave_gen_inst/_1802_ ;
 wire net137;
 wire net136;
 wire \wave_gen_inst/_1805_ ;
 wire net135;
 wire net134;
 wire \wave_gen_inst/_1808_ ;
 wire \wave_gen_inst/_1809_ ;
 wire \wave_gen_inst/_1810_ ;
 wire \wave_gen_inst/_1811_ ;
 wire \wave_gen_inst/_1812_ ;
 wire \wave_gen_inst/_1813_ ;
 wire \wave_gen_inst/_1814_ ;
 wire \wave_gen_inst/_1815_ ;
 wire \wave_gen_inst/_1816_ ;
 wire \wave_gen_inst/_1817_ ;
 wire \wave_gen_inst/_1818_ ;
 wire \wave_gen_inst/_1819_ ;
 wire \wave_gen_inst/_1820_ ;
 wire \wave_gen_inst/_1821_ ;
 wire net133;
 wire \wave_gen_inst/_1823_ ;
 wire \wave_gen_inst/_1824_ ;
 wire \wave_gen_inst/_1825_ ;
 wire \wave_gen_inst/_1826_ ;
 wire \wave_gen_inst/_1827_ ;
 wire \wave_gen_inst/_1828_ ;
 wire \wave_gen_inst/_1829_ ;
 wire \wave_gen_inst/_1830_ ;
 wire \wave_gen_inst/_1831_ ;
 wire \wave_gen_inst/_1832_ ;
 wire \wave_gen_inst/_1833_ ;
 wire net132;
 wire \wave_gen_inst/_1835_ ;
 wire \wave_gen_inst/_1836_ ;
 wire \wave_gen_inst/_1837_ ;
 wire \wave_gen_inst/_1838_ ;
 wire \wave_gen_inst/_1839_ ;
 wire \wave_gen_inst/_1840_ ;
 wire net131;
 wire \wave_gen_inst/_1842_ ;
 wire \wave_gen_inst/_1843_ ;
 wire net130;
 wire \wave_gen_inst/_1845_ ;
 wire \wave_gen_inst/_1846_ ;
 wire \wave_gen_inst/_1847_ ;
 wire \wave_gen_inst/_1848_ ;
 wire \wave_gen_inst/_1849_ ;
 wire \wave_gen_inst/_1850_ ;
 wire \wave_gen_inst/_1851_ ;
 wire \wave_gen_inst/_1852_ ;
 wire \wave_gen_inst/_1853_ ;
 wire \wave_gen_inst/_1854_ ;
 wire \wave_gen_inst/_1855_ ;
 wire \wave_gen_inst/_1856_ ;
 wire \wave_gen_inst/_1857_ ;
 wire \wave_gen_inst/_1858_ ;
 wire \wave_gen_inst/_1859_ ;
 wire \wave_gen_inst/_1860_ ;
 wire \wave_gen_inst/_1861_ ;
 wire \wave_gen_inst/_1862_ ;
 wire \wave_gen_inst/_1863_ ;
 wire \wave_gen_inst/_1864_ ;
 wire \wave_gen_inst/_1865_ ;
 wire net129;
 wire \wave_gen_inst/_1867_ ;
 wire \wave_gen_inst/_1868_ ;
 wire \wave_gen_inst/_1869_ ;
 wire \wave_gen_inst/_1870_ ;
 wire \wave_gen_inst/_1871_ ;
 wire \wave_gen_inst/_1872_ ;
 wire \wave_gen_inst/_1873_ ;
 wire \wave_gen_inst/_1874_ ;
 wire \wave_gen_inst/_1875_ ;
 wire \wave_gen_inst/_1876_ ;
 wire \wave_gen_inst/_1877_ ;
 wire \wave_gen_inst/_1878_ ;
 wire \wave_gen_inst/_1879_ ;
 wire \wave_gen_inst/_1880_ ;
 wire \wave_gen_inst/_1881_ ;
 wire \wave_gen_inst/_1882_ ;
 wire \wave_gen_inst/_1883_ ;
 wire \wave_gen_inst/_1884_ ;
 wire \wave_gen_inst/_1885_ ;
 wire \wave_gen_inst/_1886_ ;
 wire \wave_gen_inst/_1887_ ;
 wire \wave_gen_inst/_1888_ ;
 wire \wave_gen_inst/_1889_ ;
 wire \wave_gen_inst/_1890_ ;
 wire \wave_gen_inst/_1891_ ;
 wire \wave_gen_inst/_1892_ ;
 wire \wave_gen_inst/_1893_ ;
 wire \wave_gen_inst/_1894_ ;
 wire \wave_gen_inst/_1895_ ;
 wire \wave_gen_inst/_1896_ ;
 wire \wave_gen_inst/_1897_ ;
 wire \wave_gen_inst/_1898_ ;
 wire \wave_gen_inst/_1899_ ;
 wire \wave_gen_inst/_1900_ ;
 wire \wave_gen_inst/_1901_ ;
 wire \wave_gen_inst/_1902_ ;
 wire \wave_gen_inst/_1903_ ;
 wire \wave_gen_inst/_1904_ ;
 wire net128;
 wire \wave_gen_inst/_1906_ ;
 wire \wave_gen_inst/_1907_ ;
 wire \wave_gen_inst/_1908_ ;
 wire \wave_gen_inst/_1909_ ;
 wire net127;
 wire \wave_gen_inst/_1911_ ;
 wire \wave_gen_inst/_1912_ ;
 wire net126;
 wire net125;
 wire \wave_gen_inst/_1915_ ;
 wire \wave_gen_inst/_1916_ ;
 wire \wave_gen_inst/_1917_ ;
 wire net124;
 wire \wave_gen_inst/_1919_ ;
 wire \wave_gen_inst/_1920_ ;
 wire \wave_gen_inst/_1921_ ;
 wire \wave_gen_inst/_1922_ ;
 wire \wave_gen_inst/_1923_ ;
 wire \wave_gen_inst/_1924_ ;
 wire net123;
 wire \wave_gen_inst/_1926_ ;
 wire \wave_gen_inst/_1927_ ;
 wire \wave_gen_inst/_1928_ ;
 wire \wave_gen_inst/_1929_ ;
 wire \wave_gen_inst/_1930_ ;
 wire \wave_gen_inst/_1931_ ;
 wire \wave_gen_inst/_1932_ ;
 wire \wave_gen_inst/_1933_ ;
 wire \wave_gen_inst/_1934_ ;
 wire net122;
 wire \wave_gen_inst/_1936_ ;
 wire \wave_gen_inst/_1937_ ;
 wire \wave_gen_inst/_1938_ ;
 wire \wave_gen_inst/_1939_ ;
 wire \wave_gen_inst/_1940_ ;
 wire \wave_gen_inst/_1941_ ;
 wire \wave_gen_inst/_1942_ ;
 wire \wave_gen_inst/_1943_ ;
 wire net121;
 wire \wave_gen_inst/_1945_ ;
 wire \wave_gen_inst/_1946_ ;
 wire net120;
 wire \wave_gen_inst/_1948_ ;
 wire \wave_gen_inst/_1949_ ;
 wire \wave_gen_inst/_1950_ ;
 wire \wave_gen_inst/_1951_ ;
 wire net119;
 wire \wave_gen_inst/_1953_ ;
 wire \wave_gen_inst/_1954_ ;
 wire \wave_gen_inst/_1955_ ;
 wire \wave_gen_inst/_1956_ ;
 wire \wave_gen_inst/_1957_ ;
 wire \wave_gen_inst/_1958_ ;
 wire \wave_gen_inst/_1959_ ;
 wire \wave_gen_inst/_1960_ ;
 wire \wave_gen_inst/_1961_ ;
 wire \wave_gen_inst/_1962_ ;
 wire \wave_gen_inst/_1963_ ;
 wire \wave_gen_inst/_1964_ ;
 wire \wave_gen_inst/_1965_ ;
 wire \wave_gen_inst/_1966_ ;
 wire \wave_gen_inst/_1967_ ;
 wire \wave_gen_inst/_1968_ ;
 wire \wave_gen_inst/_1969_ ;
 wire \wave_gen_inst/_1970_ ;
 wire \wave_gen_inst/_1971_ ;
 wire \wave_gen_inst/_1972_ ;
 wire \wave_gen_inst/_1973_ ;
 wire \wave_gen_inst/_1974_ ;
 wire \wave_gen_inst/_1975_ ;
 wire \wave_gen_inst/_1976_ ;
 wire \wave_gen_inst/_1977_ ;
 wire \wave_gen_inst/_1978_ ;
 wire \wave_gen_inst/_1979_ ;
 wire \wave_gen_inst/_1980_ ;
 wire \wave_gen_inst/_1981_ ;
 wire \wave_gen_inst/_1982_ ;
 wire \wave_gen_inst/_1983_ ;
 wire \wave_gen_inst/_1984_ ;
 wire \wave_gen_inst/_1985_ ;
 wire \wave_gen_inst/_1986_ ;
 wire \wave_gen_inst/_1987_ ;
 wire \wave_gen_inst/_1988_ ;
 wire \wave_gen_inst/_1989_ ;
 wire \wave_gen_inst/_1990_ ;
 wire \wave_gen_inst/_1991_ ;
 wire \wave_gen_inst/_1992_ ;
 wire \wave_gen_inst/_1993_ ;
 wire \wave_gen_inst/_1994_ ;
 wire \wave_gen_inst/_1995_ ;
 wire \wave_gen_inst/_1996_ ;
 wire \wave_gen_inst/_1997_ ;
 wire \wave_gen_inst/_1998_ ;
 wire \wave_gen_inst/_1999_ ;
 wire \wave_gen_inst/_2000_ ;
 wire \wave_gen_inst/_2001_ ;
 wire \wave_gen_inst/_2002_ ;
 wire \wave_gen_inst/_2003_ ;
 wire \wave_gen_inst/_2004_ ;
 wire \wave_gen_inst/_2005_ ;
 wire \wave_gen_inst/_2006_ ;
 wire \wave_gen_inst/_2007_ ;
 wire \wave_gen_inst/_2008_ ;
 wire \wave_gen_inst/_2009_ ;
 wire \wave_gen_inst/_2010_ ;
 wire \wave_gen_inst/_2011_ ;
 wire \wave_gen_inst/_2012_ ;
 wire \wave_gen_inst/_2013_ ;
 wire \wave_gen_inst/_2014_ ;
 wire \wave_gen_inst/_2015_ ;
 wire \wave_gen_inst/_2016_ ;
 wire \wave_gen_inst/_2017_ ;
 wire \wave_gen_inst/_2018_ ;
 wire \wave_gen_inst/_2019_ ;
 wire \wave_gen_inst/_2020_ ;
 wire \wave_gen_inst/_2021_ ;
 wire \wave_gen_inst/_2022_ ;
 wire \wave_gen_inst/_2023_ ;
 wire \wave_gen_inst/_2024_ ;
 wire \wave_gen_inst/_2025_ ;
 wire \wave_gen_inst/_2026_ ;
 wire \wave_gen_inst/_2027_ ;
 wire \wave_gen_inst/_2028_ ;
 wire \wave_gen_inst/_2029_ ;
 wire \wave_gen_inst/_2030_ ;
 wire \wave_gen_inst/_2031_ ;
 wire \wave_gen_inst/_2032_ ;
 wire \wave_gen_inst/_2033_ ;
 wire \wave_gen_inst/_2034_ ;
 wire \wave_gen_inst/_2035_ ;
 wire \wave_gen_inst/_2036_ ;
 wire \wave_gen_inst/_2037_ ;
 wire \wave_gen_inst/_2038_ ;
 wire \wave_gen_inst/_2039_ ;
 wire \wave_gen_inst/_2040_ ;
 wire \wave_gen_inst/_2041_ ;
 wire \wave_gen_inst/_2042_ ;
 wire \wave_gen_inst/_2043_ ;
 wire \wave_gen_inst/_2044_ ;
 wire \wave_gen_inst/_2045_ ;
 wire \wave_gen_inst/_2046_ ;
 wire \wave_gen_inst/_2047_ ;
 wire \wave_gen_inst/_2048_ ;
 wire \wave_gen_inst/_2049_ ;
 wire \wave_gen_inst/_2050_ ;
 wire \wave_gen_inst/_2051_ ;
 wire \wave_gen_inst/_2052_ ;
 wire \wave_gen_inst/_2053_ ;
 wire \wave_gen_inst/_2054_ ;
 wire \wave_gen_inst/_2055_ ;
 wire \wave_gen_inst/_2056_ ;
 wire \wave_gen_inst/_2057_ ;
 wire \wave_gen_inst/_2058_ ;
 wire \wave_gen_inst/_2059_ ;
 wire \wave_gen_inst/_2060_ ;
 wire \wave_gen_inst/_2061_ ;
 wire \wave_gen_inst/_2062_ ;
 wire \wave_gen_inst/_2063_ ;
 wire \wave_gen_inst/_2064_ ;
 wire \wave_gen_inst/_2065_ ;
 wire \wave_gen_inst/_2066_ ;
 wire \wave_gen_inst/_2067_ ;
 wire \wave_gen_inst/_2068_ ;
 wire \wave_gen_inst/_2069_ ;
 wire \wave_gen_inst/_2070_ ;
 wire \wave_gen_inst/_2071_ ;
 wire \wave_gen_inst/_2072_ ;
 wire \wave_gen_inst/_2073_ ;
 wire \wave_gen_inst/_2074_ ;
 wire \wave_gen_inst/_2075_ ;
 wire \wave_gen_inst/_2076_ ;
 wire \wave_gen_inst/_2077_ ;
 wire \wave_gen_inst/_2078_ ;
 wire \wave_gen_inst/_2079_ ;
 wire \wave_gen_inst/_2080_ ;
 wire \wave_gen_inst/_2081_ ;
 wire \wave_gen_inst/_2082_ ;
 wire \wave_gen_inst/_2083_ ;
 wire \wave_gen_inst/_2084_ ;
 wire \wave_gen_inst/_2085_ ;
 wire \wave_gen_inst/_2086_ ;
 wire \wave_gen_inst/_2087_ ;
 wire \wave_gen_inst/_2088_ ;
 wire \wave_gen_inst/_2089_ ;
 wire \wave_gen_inst/_2090_ ;
 wire \wave_gen_inst/_2091_ ;
 wire \wave_gen_inst/_2092_ ;
 wire \wave_gen_inst/_2093_ ;
 wire \wave_gen_inst/_2094_ ;
 wire \wave_gen_inst/_2095_ ;
 wire \wave_gen_inst/_2096_ ;
 wire \wave_gen_inst/_2097_ ;
 wire \wave_gen_inst/_2098_ ;
 wire \wave_gen_inst/_2099_ ;
 wire \wave_gen_inst/_2100_ ;
 wire \wave_gen_inst/_2101_ ;
 wire \wave_gen_inst/_2102_ ;
 wire \wave_gen_inst/_2103_ ;
 wire \wave_gen_inst/_2104_ ;
 wire \wave_gen_inst/_2105_ ;
 wire \wave_gen_inst/_2106_ ;
 wire \wave_gen_inst/_2107_ ;
 wire \wave_gen_inst/_2108_ ;
 wire \wave_gen_inst/_2109_ ;
 wire \wave_gen_inst/_2110_ ;
 wire \wave_gen_inst/_2111_ ;
 wire \wave_gen_inst/_2112_ ;
 wire \wave_gen_inst/_2113_ ;
 wire \wave_gen_inst/_2114_ ;
 wire \wave_gen_inst/_2115_ ;
 wire \wave_gen_inst/_2116_ ;
 wire \wave_gen_inst/_2117_ ;
 wire \wave_gen_inst/_2118_ ;
 wire \wave_gen_inst/_2119_ ;
 wire \wave_gen_inst/_2120_ ;
 wire \wave_gen_inst/_2121_ ;
 wire \wave_gen_inst/_2122_ ;
 wire \wave_gen_inst/_2123_ ;
 wire \wave_gen_inst/_2124_ ;
 wire \wave_gen_inst/_2125_ ;
 wire \wave_gen_inst/_2126_ ;
 wire \wave_gen_inst/_2127_ ;
 wire \wave_gen_inst/_2128_ ;
 wire \wave_gen_inst/_2129_ ;
 wire \wave_gen_inst/_2130_ ;
 wire \wave_gen_inst/_2131_ ;
 wire \wave_gen_inst/_2132_ ;
 wire \wave_gen_inst/_2133_ ;
 wire \wave_gen_inst/_2134_ ;
 wire \wave_gen_inst/_2135_ ;
 wire \wave_gen_inst/_2136_ ;
 wire \wave_gen_inst/_2137_ ;
 wire \wave_gen_inst/_2138_ ;
 wire \wave_gen_inst/_2139_ ;
 wire \wave_gen_inst/_2140_ ;
 wire \wave_gen_inst/_2141_ ;
 wire \wave_gen_inst/_2142_ ;
 wire \wave_gen_inst/_2143_ ;
 wire \wave_gen_inst/_2144_ ;
 wire \wave_gen_inst/_2145_ ;
 wire \wave_gen_inst/_2146_ ;
 wire \wave_gen_inst/_2147_ ;
 wire \wave_gen_inst/_2148_ ;
 wire \wave_gen_inst/_2149_ ;
 wire \wave_gen_inst/_2150_ ;
 wire \wave_gen_inst/_2151_ ;
 wire \wave_gen_inst/_2152_ ;
 wire \wave_gen_inst/_2153_ ;
 wire \wave_gen_inst/_2154_ ;
 wire \wave_gen_inst/_2155_ ;
 wire \wave_gen_inst/_2156_ ;
 wire \wave_gen_inst/_2157_ ;
 wire \wave_gen_inst/_2158_ ;
 wire \wave_gen_inst/_2159_ ;
 wire \wave_gen_inst/_2160_ ;
 wire \wave_gen_inst/_2161_ ;
 wire \wave_gen_inst/_2162_ ;
 wire \wave_gen_inst/_2163_ ;
 wire \wave_gen_inst/_2164_ ;
 wire \wave_gen_inst/_2165_ ;
 wire \wave_gen_inst/_2166_ ;
 wire \wave_gen_inst/_2167_ ;
 wire \wave_gen_inst/_2168_ ;
 wire \wave_gen_inst/_2169_ ;
 wire \wave_gen_inst/_2170_ ;
 wire \wave_gen_inst/_2171_ ;
 wire \wave_gen_inst/_2172_ ;
 wire \wave_gen_inst/_2173_ ;
 wire \wave_gen_inst/_2174_ ;
 wire \wave_gen_inst/_2175_ ;
 wire \wave_gen_inst/_2176_ ;
 wire \wave_gen_inst/_2177_ ;
 wire \wave_gen_inst/_2178_ ;
 wire \wave_gen_inst/_2179_ ;
 wire \wave_gen_inst/_2180_ ;
 wire \wave_gen_inst/_2181_ ;
 wire \wave_gen_inst/_2182_ ;
 wire \wave_gen_inst/_2183_ ;
 wire \wave_gen_inst/_2184_ ;
 wire \wave_gen_inst/_2185_ ;
 wire \wave_gen_inst/_2186_ ;
 wire \wave_gen_inst/_2187_ ;
 wire \wave_gen_inst/_2188_ ;
 wire \wave_gen_inst/_2189_ ;
 wire \wave_gen_inst/_2190_ ;
 wire \wave_gen_inst/_2191_ ;
 wire \wave_gen_inst/_2192_ ;
 wire \wave_gen_inst/_2193_ ;
 wire \wave_gen_inst/_2194_ ;
 wire \wave_gen_inst/_2195_ ;
 wire net118;
 wire net117;
 wire net116;
 wire net115;
 wire net114;
 wire net113;
 wire net112;
 wire net473;
 wire \wave_gen_inst/changed ;
 wire \wave_gen_inst/counter[0] ;
 wire \wave_gen_inst/counter[10] ;
 wire \wave_gen_inst/counter[11] ;
 wire \wave_gen_inst/counter[12] ;
 wire \wave_gen_inst/counter[13] ;
 wire \wave_gen_inst/counter[14] ;
 wire \wave_gen_inst/counter[15] ;
 wire \wave_gen_inst/counter[16] ;
 wire \wave_gen_inst/counter[17] ;
 wire \wave_gen_inst/counter[18] ;
 wire \wave_gen_inst/counter[19] ;
 wire \wave_gen_inst/counter[1] ;
 wire \wave_gen_inst/counter[20] ;
 wire \wave_gen_inst/counter[21] ;
 wire \wave_gen_inst/counter[22] ;
 wire \wave_gen_inst/counter[23] ;
 wire \wave_gen_inst/counter[24] ;
 wire \wave_gen_inst/counter[25] ;
 wire \wave_gen_inst/counter[26] ;
 wire \wave_gen_inst/counter[27] ;
 wire \wave_gen_inst/counter[28] ;
 wire \wave_gen_inst/counter[29] ;
 wire \wave_gen_inst/counter[2] ;
 wire \wave_gen_inst/counter[30] ;
 wire \wave_gen_inst/counter[31] ;
 wire \wave_gen_inst/counter[3] ;
 wire \wave_gen_inst/counter[4] ;
 wire \wave_gen_inst/counter[5] ;
 wire \wave_gen_inst/counter[6] ;
 wire \wave_gen_inst/counter[7] ;
 wire \wave_gen_inst/counter[8] ;
 wire \wave_gen_inst/counter[9] ;
 wire \wave_gen_inst/param1[0] ;
 wire \wave_gen_inst/param1[10] ;
 wire \wave_gen_inst/param1[11] ;
 wire \wave_gen_inst/param1[1] ;
 wire \wave_gen_inst/param1[2] ;
 wire \wave_gen_inst/param1[3] ;
 wire \wave_gen_inst/param1[4] ;
 wire \wave_gen_inst/param1[5] ;
 wire \wave_gen_inst/param1[6] ;
 wire \wave_gen_inst/param1[7] ;
 wire \wave_gen_inst/param1[8] ;
 wire \wave_gen_inst/param1[9] ;
 wire \wave_gen_inst/param2[0] ;
 wire \wave_gen_inst/param2[10] ;
 wire \wave_gen_inst/param2[11] ;
 wire \wave_gen_inst/param2[1] ;
 wire \wave_gen_inst/param2[2] ;
 wire \wave_gen_inst/param2[3] ;
 wire \wave_gen_inst/param2[4] ;
 wire \wave_gen_inst/param2[5] ;
 wire \wave_gen_inst/param2[6] ;
 wire \wave_gen_inst/param2[7] ;
 wire \wave_gen_inst/param2[8] ;
 wire \wave_gen_inst/param2[9] ;
 wire \wave_gen_inst/pp ;
 wire \wave_gen_inst/rom_output[0] ;
 wire \wave_gen_inst/rom_output[10] ;
 wire \wave_gen_inst/rom_output[1] ;
 wire \wave_gen_inst/rom_output[2] ;
 wire \wave_gen_inst/rom_output[3] ;
 wire \wave_gen_inst/rom_output[4] ;
 wire \wave_gen_inst/rom_output[5] ;
 wire \wave_gen_inst/rom_output[6] ;
 wire \wave_gen_inst/rom_output[7] ;
 wire \wave_gen_inst/rom_output[8] ;
 wire \wave_gen_inst/rom_output[9] ;
 wire \wave_gen_inst/sign ;
 wire \wave_gen_inst/sine_phase[0] ;
 wire \wave_gen_inst/sine_phase[1] ;
 wire \wave_gen_inst/sine_phase[2] ;
 wire \wave_gen_inst/sine_phase[3] ;
 wire \wave_gen_inst/sine_phase[4] ;
 wire \wave_gen_inst/sine_phase[5] ;
 wire \wave_gen_inst/sine_phase[6] ;
 wire \wave_gen_inst/rom/_000_ ;
 wire \wave_gen_inst/rom/_001_ ;
 wire \wave_gen_inst/rom/_002_ ;
 wire \wave_gen_inst/rom/_003_ ;
 wire \wave_gen_inst/rom/_004_ ;
 wire \wave_gen_inst/rom/_005_ ;
 wire \wave_gen_inst/rom/_006_ ;
 wire \wave_gen_inst/rom/_007_ ;
 wire \wave_gen_inst/rom/_008_ ;
 wire \wave_gen_inst/rom/_009_ ;
 wire net2;
 wire \wave_gen_inst/rom/_011_ ;
 wire \wave_gen_inst/rom/_012_ ;
 wire \wave_gen_inst/rom/_013_ ;
 wire \wave_gen_inst/rom/_014_ ;
 wire \wave_gen_inst/rom/_015_ ;
 wire \wave_gen_inst/rom/_016_ ;
 wire \wave_gen_inst/rom/_017_ ;
 wire \wave_gen_inst/rom/_018_ ;
 wire \wave_gen_inst/rom/_019_ ;
 wire net1;
 wire \wave_gen_inst/rom/_021_ ;
 wire \wave_gen_inst/rom/_022_ ;
 wire \wave_gen_inst/rom/_023_ ;
 wire \wave_gen_inst/rom/_024_ ;
 wire \wave_gen_inst/rom/_025_ ;
 wire \wave_gen_inst/rom/_026_ ;
 wire \wave_gen_inst/rom/_027_ ;
 wire \wave_gen_inst/rom/_029_ ;
 wire \wave_gen_inst/rom/_030_ ;
 wire \wave_gen_inst/rom/_031_ ;
 wire \wave_gen_inst/rom/_032_ ;
 wire \wave_gen_inst/rom/_033_ ;
 wire \wave_gen_inst/rom/_034_ ;
 wire \wave_gen_inst/rom/_035_ ;
 wire \wave_gen_inst/rom/_036_ ;
 wire \wave_gen_inst/rom/_037_ ;
 wire \wave_gen_inst/rom/_038_ ;
 wire \wave_gen_inst/rom/_039_ ;
 wire \wave_gen_inst/rom/_040_ ;
 wire \wave_gen_inst/rom/_041_ ;
 wire \wave_gen_inst/rom/_042_ ;
 wire \wave_gen_inst/rom/_043_ ;
 wire \wave_gen_inst/rom/_044_ ;
 wire \wave_gen_inst/rom/_045_ ;
 wire \wave_gen_inst/rom/_046_ ;
 wire \wave_gen_inst/rom/_047_ ;
 wire \wave_gen_inst/rom/_048_ ;
 wire \wave_gen_inst/rom/_049_ ;
 wire \wave_gen_inst/rom/_050_ ;
 wire \wave_gen_inst/rom/_051_ ;
 wire \wave_gen_inst/rom/_052_ ;
 wire \wave_gen_inst/rom/_053_ ;
 wire \wave_gen_inst/rom/_054_ ;
 wire \wave_gen_inst/rom/_055_ ;
 wire \wave_gen_inst/rom/_056_ ;
 wire \wave_gen_inst/rom/_057_ ;
 wire \wave_gen_inst/rom/_058_ ;
 wire \wave_gen_inst/rom/_059_ ;
 wire \wave_gen_inst/rom/_060_ ;
 wire \wave_gen_inst/rom/_061_ ;
 wire \wave_gen_inst/rom/_062_ ;
 wire \wave_gen_inst/rom/_063_ ;
 wire \wave_gen_inst/rom/_064_ ;
 wire \wave_gen_inst/rom/_065_ ;
 wire \wave_gen_inst/rom/_066_ ;
 wire \wave_gen_inst/rom/_067_ ;
 wire \wave_gen_inst/rom/_068_ ;
 wire \wave_gen_inst/rom/_069_ ;
 wire \wave_gen_inst/rom/_070_ ;
 wire \wave_gen_inst/rom/_071_ ;
 wire \wave_gen_inst/rom/_072_ ;
 wire \wave_gen_inst/rom/_073_ ;
 wire \wave_gen_inst/rom/_074_ ;
 wire \wave_gen_inst/rom/_075_ ;
 wire \wave_gen_inst/rom/_076_ ;
 wire \wave_gen_inst/rom/_077_ ;
 wire \wave_gen_inst/rom/_078_ ;
 wire \wave_gen_inst/rom/_079_ ;
 wire \wave_gen_inst/rom/_080_ ;
 wire \wave_gen_inst/rom/_081_ ;
 wire \wave_gen_inst/rom/_082_ ;
 wire \wave_gen_inst/rom/_083_ ;
 wire \wave_gen_inst/rom/_084_ ;
 wire \wave_gen_inst/rom/_085_ ;
 wire \wave_gen_inst/rom/_086_ ;
 wire \wave_gen_inst/rom/_087_ ;
 wire \wave_gen_inst/rom/_088_ ;
 wire \wave_gen_inst/rom/_089_ ;
 wire \wave_gen_inst/rom/_090_ ;
 wire \wave_gen_inst/rom/_091_ ;
 wire \wave_gen_inst/rom/_092_ ;
 wire \wave_gen_inst/rom/_093_ ;
 wire \wave_gen_inst/rom/_094_ ;
 wire \wave_gen_inst/rom/_095_ ;
 wire net28;
 wire \wave_gen_inst/rom/_097_ ;
 wire \wave_gen_inst/rom/_098_ ;
 wire \wave_gen_inst/rom/_099_ ;
 wire \wave_gen_inst/rom/_100_ ;
 wire \wave_gen_inst/rom/_101_ ;
 wire \wave_gen_inst/rom/_102_ ;
 wire \wave_gen_inst/rom/_103_ ;
 wire \wave_gen_inst/rom/_104_ ;
 wire \wave_gen_inst/rom/_105_ ;
 wire \wave_gen_inst/rom/_106_ ;
 wire net27;
 wire \wave_gen_inst/rom/_108_ ;
 wire \wave_gen_inst/rom/_109_ ;
 wire \wave_gen_inst/rom/_110_ ;
 wire \wave_gen_inst/rom/_111_ ;
 wire \wave_gen_inst/rom/_112_ ;
 wire \wave_gen_inst/rom/_113_ ;
 wire \wave_gen_inst/rom/_114_ ;
 wire \wave_gen_inst/rom/_115_ ;
 wire \wave_gen_inst/rom/_116_ ;
 wire net26;
 wire \wave_gen_inst/rom/_118_ ;
 wire \wave_gen_inst/rom/_119_ ;
 wire \wave_gen_inst/rom/_120_ ;
 wire \wave_gen_inst/rom/_121_ ;
 wire \wave_gen_inst/rom/_122_ ;
 wire \wave_gen_inst/rom/_123_ ;
 wire \wave_gen_inst/rom/_124_ ;
 wire \wave_gen_inst/rom/_125_ ;
 wire \wave_gen_inst/rom/_126_ ;
 wire \wave_gen_inst/rom/_127_ ;
 wire net25;
 wire \wave_gen_inst/rom/_129_ ;
 wire \wave_gen_inst/rom/_130_ ;
 wire \wave_gen_inst/rom/_131_ ;
 wire \wave_gen_inst/rom/_132_ ;
 wire \wave_gen_inst/rom/_133_ ;
 wire \wave_gen_inst/rom/_134_ ;
 wire \wave_gen_inst/rom/_135_ ;
 wire \wave_gen_inst/rom/_136_ ;
 wire \wave_gen_inst/rom/_137_ ;
 wire net24;
 wire \wave_gen_inst/rom/_139_ ;
 wire \wave_gen_inst/rom/_140_ ;
 wire \wave_gen_inst/rom/_141_ ;
 wire \wave_gen_inst/rom/_142_ ;
 wire \wave_gen_inst/rom/_143_ ;
 wire \wave_gen_inst/rom/_144_ ;
 wire \wave_gen_inst/rom/_145_ ;
 wire \wave_gen_inst/rom/_146_ ;
 wire \wave_gen_inst/rom/_147_ ;
 wire net23;
 wire \wave_gen_inst/rom/_149_ ;
 wire \wave_gen_inst/rom/_150_ ;
 wire \wave_gen_inst/rom/_151_ ;
 wire \wave_gen_inst/rom/_152_ ;
 wire \wave_gen_inst/rom/_153_ ;
 wire \wave_gen_inst/rom/_154_ ;
 wire \wave_gen_inst/rom/_155_ ;
 wire \wave_gen_inst/rom/_156_ ;
 wire \wave_gen_inst/rom/_157_ ;
 wire net22;
 wire \wave_gen_inst/rom/_159_ ;
 wire \wave_gen_inst/rom/_160_ ;
 wire \wave_gen_inst/rom/_161_ ;
 wire \wave_gen_inst/rom/_162_ ;
 wire \wave_gen_inst/rom/_163_ ;
 wire \wave_gen_inst/rom/_164_ ;
 wire net21;
 wire \wave_gen_inst/rom/_166_ ;
 wire net20;
 wire net19;
 wire \wave_gen_inst/rom/_169_ ;
 wire net18;
 wire \wave_gen_inst/rom/_171_ ;
 wire net17;
 wire net16;
 wire net15;
 wire \wave_gen_inst/rom/_175_ ;
 wire net14;
 wire net13;
 wire \wave_gen_inst/rom/_178_ ;
 wire \wave_gen_inst/rom/_179_ ;
 wire \wave_gen_inst/rom/_180_ ;
 wire \wave_gen_inst/rom/_181_ ;
 wire \wave_gen_inst/rom/_182_ ;
 wire net12;
 wire \wave_gen_inst/rom/_184_ ;
 wire \wave_gen_inst/rom/_185_ ;
 wire \wave_gen_inst/rom/_186_ ;
 wire \wave_gen_inst/rom/_187_ ;
 wire net11;
 wire \wave_gen_inst/rom/_189_ ;
 wire \wave_gen_inst/rom/_190_ ;
 wire \wave_gen_inst/rom/_191_ ;
 wire \wave_gen_inst/rom/_192_ ;
 wire \wave_gen_inst/rom/_193_ ;
 wire \wave_gen_inst/rom/_194_ ;
 wire \wave_gen_inst/rom/_195_ ;
 wire \wave_gen_inst/rom/_196_ ;
 wire net10;
 wire \wave_gen_inst/rom/_198_ ;
 wire \wave_gen_inst/rom/_199_ ;
 wire \wave_gen_inst/rom/_200_ ;
 wire \wave_gen_inst/rom/_201_ ;
 wire net9;
 wire \wave_gen_inst/rom/_203_ ;
 wire net8;
 wire \wave_gen_inst/rom/_205_ ;
 wire net7;
 wire \wave_gen_inst/rom/_207_ ;
 wire \wave_gen_inst/rom/_208_ ;
 wire \wave_gen_inst/rom/_209_ ;
 wire \wave_gen_inst/rom/_210_ ;
 wire \wave_gen_inst/rom/_211_ ;
 wire \wave_gen_inst/rom/_212_ ;
 wire net6;
 wire \wave_gen_inst/rom/_214_ ;
 wire \wave_gen_inst/rom/_215_ ;
 wire \wave_gen_inst/rom/_216_ ;
 wire net5;
 wire \wave_gen_inst/rom/_218_ ;
 wire \wave_gen_inst/rom/_219_ ;
 wire \wave_gen_inst/rom/_220_ ;
 wire \wave_gen_inst/rom/_221_ ;
 wire \wave_gen_inst/rom/_222_ ;
 wire net4;
 wire \wave_gen_inst/rom/_224_ ;
 wire net3;
 wire \wave_gen_inst/rom/_226_ ;
 wire \wave_gen_inst/rom/_227_ ;
 wire \wave_gen_inst/rom/_228_ ;
 wire \wave_gen_inst/rom/_229_ ;
 wire \wave_gen_inst/rom/_230_ ;
 wire \wave_gen_inst/rom/_231_ ;
 wire \wave_gen_inst/rom/_232_ ;
 wire \wave_gen_inst/rom/_233_ ;
 wire \wave_gen_inst/rom/_234_ ;
 wire \wave_gen_inst/rom/_235_ ;
 wire \wave_gen_inst/rom/_236_ ;
 wire \wave_gen_inst/rom/_237_ ;
 wire net488;
 wire [31:0] \soc/cpu/eoi ;
 wire [31:0] \soc/cpu/mem_la_addr ;
 wire [31:0] \soc/cpu/mem_la_wdata ;
 wire [3:0] \soc/cpu/mem_la_wstrb ;
 wire [31:0] \soc/cpu/pcpi_rs1 ;
 wire [31:0] \soc/cpu/pcpi_rs2 ;

 sky130_fd_sc_hd__nand2_1 _198_ (.A(net944),
    .B(\reset_cnt[0] ),
    .Y(_071_));
 sky130_fd_sc_hd__nand4_1 _199_ (.A(\reset_cnt[3] ),
    .B(\reset_cnt[2] ),
    .C(\reset_cnt[5] ),
    .D(\reset_cnt[4] ),
    .Y(_072_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _200_ (.A(_071_),
    .SLEEP(_072_),
    .X(_073_));
 sky130_fd_sc_hd__clkinv_16 _201_ (.A(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__clkinv_4 _203_ (.A(\gpio[6] ),
    .Y(net10));
 sky130_fd_sc_hd__inv_4 _204_ (.A(\gpio[7] ),
    .Y(net9));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 _205_ (.A(_072_),
    .SLEEP(_071_),
    .X(_075_));
 sky130_fd_sc_hd__nor2_1 _206_ (.A(\reset_cnt[1] ),
    .B(\reset_cnt[0] ),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_1 _207_ (.A(_075_),
    .B(_076_),
    .Y(_001_));
 sky130_fd_sc_hd__xor2_1 _208_ (.A(\reset_cnt[2] ),
    .B(_075_),
    .X(_002_));
 sky130_fd_sc_hd__a21oi_1 _209_ (.A1(\reset_cnt[2] ),
    .A2(_075_),
    .B1(\reset_cnt[3] ),
    .Y(_077_));
 sky130_fd_sc_hd__nand3_1 _210_ (.A(net837),
    .B(\reset_cnt[2] ),
    .C(_075_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2b_1 _211_ (.A(_077_),
    .B_N(_078_),
    .Y(_003_));
 sky130_fd_sc_hd__xnor2_1 _212_ (.A(\reset_cnt[4] ),
    .B(net838),
    .Y(_004_));
 sky130_fd_sc_hd__a41o_1 _213_ (.A1(\reset_cnt[3] ),
    .A2(\reset_cnt[2] ),
    .A3(\reset_cnt[4] ),
    .A4(_075_),
    .B1(\reset_cnt[5] ),
    .X(_005_));
 sky130_fd_sc_hd__nand2_1 _214_ (.A(\reset_cnt[0] ),
    .B(_073_),
    .Y(_000_));
 sky130_fd_sc_hd__nor4_4 _215_ (.A(net739),
    .B(\iomem_addr[28] ),
    .C(\iomem_addr[31] ),
    .D(net717),
    .Y(_079_));
 sky130_fd_sc_hd__nor2_1 _216_ (.A(\iomem_addr[24] ),
    .B(net701),
    .Y(_080_));
 sky130_fd_sc_hd__nand4b_4 _217_ (.A_N(net492),
    .B(net809),
    .C(net718),
    .D(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__mux2_1 _219_ (.A0(net15),
    .A1(\gpio[0] ),
    .S(_081_),
    .X(_083_));
 sky130_fd_sc_hd__nor4bb_4 _220_ (.A(net701),
    .B(net941),
    .C_N(net492),
    .D_N(\iomem_addr[24] ),
    .Y(_084_));
 sky130_fd_sc_hd__nand2_1 _221_ (.A(net718),
    .B(net702),
    .Y(_085_));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 _222_ (.A(iomem_valid),
    .SLEEP(net808),
    .X(_086_));
 sky130_fd_sc_hd__inv_1 _223_ (.A(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a211oi_4 _224_ (.A1(_085_),
    .A2(_081_),
    .B1(_087_),
    .C1(_073_),
    .Y(_088_));
 sky130_fd_sc_hd__mux2_1 _226_ (.A0(\iomem_rdata[0] ),
    .A1(_083_),
    .S(net120),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _227_ (.A0(net768),
    .A1(net4),
    .S(net151),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _228_ (.A0(\iomem_rdata[1] ),
    .A1(net769),
    .S(net121),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _229_ (.A0(net757),
    .A1(net5),
    .S(net151),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _230_ (.A0(\iomem_rdata[2] ),
    .A1(net758),
    .S(net122),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _231_ (.A0(net40),
    .A1(net6),
    .S(net151),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _232_ (.A0(\iomem_rdata[3] ),
    .A1(_092_),
    .S(net122),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _233_ (.A0(net41),
    .A1(net7),
    .S(_081_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _234_ (.A0(\iomem_rdata[4] ),
    .A1(_093_),
    .S(net120),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _235_ (.A0(net42),
    .A1(net8),
    .S(_081_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _236_ (.A0(\iomem_rdata[5] ),
    .A1(_094_),
    .S(net120),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _237_ (.A0(net796),
    .A1(\gpio[6] ),
    .S(net151),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _238_ (.A0(\iomem_rdata[6] ),
    .A1(net797),
    .S(net121),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _239_ (.A0(net44),
    .A1(\gpio[7] ),
    .S(_081_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _240_ (.A0(\iomem_rdata[7] ),
    .A1(_096_),
    .S(net120),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _241_ (.A0(net45),
    .A1(\gpio[8] ),
    .S(_081_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _242_ (.A0(\iomem_rdata[8] ),
    .A1(_097_),
    .S(net120),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _243_ (.A0(net46),
    .A1(\gpio[9] ),
    .S(net151),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _245_ (.A0(\iomem_rdata[9] ),
    .A1(net810),
    .S(net122),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _247_ (.A0(net16),
    .A1(\gpio[10] ),
    .S(net151),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _248_ (.A0(\iomem_rdata[10] ),
    .A1(_101_),
    .S(net122),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _249_ (.A0(net17),
    .A1(\gpio[11] ),
    .S(_081_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _250_ (.A0(\iomem_rdata[11] ),
    .A1(_102_),
    .S(net120),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _251_ (.A0(net18),
    .A1(\gpio[12] ),
    .S(_081_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _252_ (.A0(\iomem_rdata[12] ),
    .A1(_103_),
    .S(net120),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _253_ (.A0(net19),
    .A1(\gpio[13] ),
    .S(_081_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(\iomem_rdata[13] ),
    .A1(_104_),
    .S(net120),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _255_ (.A0(net20),
    .A1(\gpio[14] ),
    .S(net151),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _256_ (.A0(\iomem_rdata[14] ),
    .A1(_105_),
    .S(net121),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _257_ (.A0(net21),
    .A1(\gpio[15] ),
    .S(_081_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(\iomem_rdata[15] ),
    .A1(_106_),
    .S(net120),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _259_ (.A0(net22),
    .A1(\gpio[16] ),
    .S(_081_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _260_ (.A0(\iomem_rdata[16] ),
    .A1(_107_),
    .S(net120),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(net23),
    .A1(\gpio[17] ),
    .S(net151),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _262_ (.A0(\iomem_rdata[17] ),
    .A1(_108_),
    .S(net121),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _263_ (.A0(net24),
    .A1(\gpio[18] ),
    .S(net151),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _264_ (.A0(\iomem_rdata[18] ),
    .A1(_109_),
    .S(net121),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _265_ (.A0(net25),
    .A1(\gpio[19] ),
    .S(net151),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _267_ (.A0(\iomem_rdata[19] ),
    .A1(_110_),
    .S(net122),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(net27),
    .A1(\gpio[20] ),
    .S(net151),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _270_ (.A0(\iomem_rdata[20] ),
    .A1(_113_),
    .S(net122),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _271_ (.A0(net28),
    .A1(\gpio[21] ),
    .S(_081_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _272_ (.A0(\iomem_rdata[21] ),
    .A1(_114_),
    .S(net120),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(net29),
    .A1(\gpio[22] ),
    .S(net151),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _274_ (.A0(\iomem_rdata[22] ),
    .A1(_115_),
    .S(net121),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(net30),
    .A1(\gpio[23] ),
    .S(_081_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _276_ (.A0(\iomem_rdata[23] ),
    .A1(_116_),
    .S(net120),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(net31),
    .A1(net869),
    .S(net151),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(\iomem_rdata[24] ),
    .A1(_117_),
    .S(_088_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(net32),
    .A1(\gpio[25] ),
    .S(net151),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _280_ (.A0(\iomem_rdata[25] ),
    .A1(_118_),
    .S(net122),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(net33),
    .A1(\gpio[26] ),
    .S(net151),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _282_ (.A0(\iomem_rdata[26] ),
    .A1(_119_),
    .S(net121),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(net34),
    .A1(\gpio[27] ),
    .S(net151),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(\iomem_rdata[27] ),
    .A1(_120_),
    .S(_088_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(net35),
    .A1(\gpio[28] ),
    .S(net151),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _286_ (.A0(\iomem_rdata[28] ),
    .A1(_121_),
    .S(_088_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(net36),
    .A1(\gpio[29] ),
    .S(_081_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(\iomem_rdata[29] ),
    .A1(_122_),
    .S(_088_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(net38),
    .A1(net704),
    .S(net151),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(\iomem_rdata[30] ),
    .A1(net705),
    .S(net121),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(net39),
    .A1(\gpio[31] ),
    .S(_081_),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(\iomem_rdata[31] ),
    .A1(_124_),
    .S(_088_),
    .X(_045_));
 sky130_fd_sc_hd__a21o_1 _293_ (.A1(iomem_ready),
    .A2(_073_),
    .B1(_088_),
    .X(_062_));
 sky130_fd_sc_hd__inv_1 _294_ (.A(\gpio[8] ),
    .Y(_125_));
 sky130_fd_sc_hd__nand4_4 _295_ (.A(net407),
    .B(net718),
    .C(net702),
    .D(_086_),
    .Y(_126_));
 sky130_fd_sc_hd__o21ai_0 _297_ (.A1(net251),
    .A2(net719),
    .B1(_074_),
    .Y(_128_));
 sky130_fd_sc_hd__a21oi_1 _298_ (.A1(_125_),
    .A2(net719),
    .B1(_128_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_1 _299_ (.A(\gpio[9] ),
    .Y(_129_));
 sky130_fd_sc_hd__o21ai_0 _300_ (.A1(net238),
    .A2(net719),
    .B1(_074_),
    .Y(_130_));
 sky130_fd_sc_hd__a21oi_1 _301_ (.A1(_129_),
    .A2(net719),
    .B1(_130_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_1 _302_ (.A(\gpio[10] ),
    .Y(_131_));
 sky130_fd_sc_hd__o21ai_0 _303_ (.A1(net235),
    .A2(net719),
    .B1(_074_),
    .Y(_132_));
 sky130_fd_sc_hd__a21oi_1 _304_ (.A1(_131_),
    .A2(net719),
    .B1(_132_),
    .Y(_008_));
 sky130_fd_sc_hd__inv_1 _305_ (.A(\gpio[11] ),
    .Y(_133_));
 sky130_fd_sc_hd__o21ai_0 _306_ (.A1(net233),
    .A2(_126_),
    .B1(_074_),
    .Y(_134_));
 sky130_fd_sc_hd__a21oi_1 _307_ (.A1(_133_),
    .A2(_126_),
    .B1(_134_),
    .Y(_009_));
 sky130_fd_sc_hd__inv_1 _308_ (.A(\gpio[12] ),
    .Y(_135_));
 sky130_fd_sc_hd__o21ai_0 _309_ (.A1(net229),
    .A2(_126_),
    .B1(_074_),
    .Y(_136_));
 sky130_fd_sc_hd__a21oi_1 _310_ (.A1(_135_),
    .A2(_126_),
    .B1(_136_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_1 _311_ (.A(\gpio[13] ),
    .Y(_137_));
 sky130_fd_sc_hd__o21ai_0 _312_ (.A1(net225),
    .A2(_126_),
    .B1(_074_),
    .Y(_138_));
 sky130_fd_sc_hd__a21oi_1 _313_ (.A1(_137_),
    .A2(_126_),
    .B1(_138_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_1 _314_ (.A(\gpio[14] ),
    .Y(_139_));
 sky130_fd_sc_hd__o21ai_0 _315_ (.A1(net220),
    .A2(net719),
    .B1(_074_),
    .Y(_140_));
 sky130_fd_sc_hd__a21oi_1 _316_ (.A1(_139_),
    .A2(net719),
    .B1(_140_),
    .Y(_012_));
 sky130_fd_sc_hd__inv_1 _317_ (.A(\gpio[15] ),
    .Y(_141_));
 sky130_fd_sc_hd__o21ai_0 _318_ (.A1(net218),
    .A2(_126_),
    .B1(_074_),
    .Y(_142_));
 sky130_fd_sc_hd__a21oi_1 _319_ (.A1(_141_),
    .A2(_126_),
    .B1(_142_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_1 _320_ (.A(\gpio[24] ),
    .Y(_143_));
 sky130_fd_sc_hd__nand4_4 _321_ (.A(net398),
    .B(_079_),
    .C(_084_),
    .D(_086_),
    .Y(_144_));
 sky130_fd_sc_hd__o21ai_0 _323_ (.A1(net185),
    .A2(_144_),
    .B1(_074_),
    .Y(_146_));
 sky130_fd_sc_hd__a21oi_1 _324_ (.A1(_143_),
    .A2(_144_),
    .B1(_146_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_1 _325_ (.A(\gpio[25] ),
    .Y(_147_));
 sky130_fd_sc_hd__o21ai_0 _327_ (.A1(net182),
    .A2(_144_),
    .B1(_074_),
    .Y(_149_));
 sky130_fd_sc_hd__a21oi_1 _328_ (.A1(_147_),
    .A2(_144_),
    .B1(_149_),
    .Y(_047_));
 sky130_fd_sc_hd__inv_1 _329_ (.A(\gpio[26] ),
    .Y(_150_));
 sky130_fd_sc_hd__o21ai_0 _330_ (.A1(net179),
    .A2(_144_),
    .B1(_074_),
    .Y(_151_));
 sky130_fd_sc_hd__a21oi_1 _331_ (.A1(_150_),
    .A2(_144_),
    .B1(_151_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_1 _332_ (.A(\gpio[27] ),
    .Y(_152_));
 sky130_fd_sc_hd__o21ai_0 _333_ (.A1(net176),
    .A2(_144_),
    .B1(_074_),
    .Y(_153_));
 sky130_fd_sc_hd__a21oi_1 _334_ (.A1(_152_),
    .A2(_144_),
    .B1(_153_),
    .Y(_049_));
 sky130_fd_sc_hd__inv_1 _335_ (.A(\gpio[28] ),
    .Y(_154_));
 sky130_fd_sc_hd__o21ai_0 _336_ (.A1(net173),
    .A2(_144_),
    .B1(_074_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_1 _337_ (.A1(_154_),
    .A2(_144_),
    .B1(_155_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_1 _338_ (.A(\gpio[29] ),
    .Y(_156_));
 sky130_fd_sc_hd__o21ai_0 _339_ (.A1(net170),
    .A2(_144_),
    .B1(_074_),
    .Y(_157_));
 sky130_fd_sc_hd__a21oi_1 _340_ (.A1(_156_),
    .A2(_144_),
    .B1(_157_),
    .Y(_051_));
 sky130_fd_sc_hd__nand4_1 _341_ (.A(net399),
    .B(_079_),
    .C(_084_),
    .D(_086_),
    .Y(_158_));
 sky130_fd_sc_hd__mux2i_1 _342_ (.A0(net167),
    .A1(\gpio[30] ),
    .S(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _343_ (.A(_073_),
    .B(_159_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_1 _344_ (.A(\gpio[31] ),
    .Y(_160_));
 sky130_fd_sc_hd__o21ai_0 _345_ (.A1(net165),
    .A2(_144_),
    .B1(_074_),
    .Y(_161_));
 sky130_fd_sc_hd__a21oi_1 _346_ (.A1(_160_),
    .A2(_144_),
    .B1(_161_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_1 _347_ (.A(\gpio[16] ),
    .Y(_162_));
 sky130_fd_sc_hd__nand4_4 _348_ (.A(net403),
    .B(_079_),
    .C(_084_),
    .D(_086_),
    .Y(_163_));
 sky130_fd_sc_hd__o21ai_0 _350_ (.A1(net214),
    .A2(_163_),
    .B1(_074_),
    .Y(_165_));
 sky130_fd_sc_hd__a21oi_1 _351_ (.A1(_162_),
    .A2(net942),
    .B1(_165_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_1 _352_ (.A(\gpio[17] ),
    .Y(_166_));
 sky130_fd_sc_hd__o21ai_0 _353_ (.A1(net209),
    .A2(_163_),
    .B1(_074_),
    .Y(_167_));
 sky130_fd_sc_hd__a21oi_1 _354_ (.A1(_166_),
    .A2(_163_),
    .B1(_167_),
    .Y(_055_));
 sky130_fd_sc_hd__inv_1 _355_ (.A(\gpio[18] ),
    .Y(_168_));
 sky130_fd_sc_hd__o21ai_0 _356_ (.A1(net206),
    .A2(_163_),
    .B1(_074_),
    .Y(_169_));
 sky130_fd_sc_hd__a21oi_1 _357_ (.A1(_168_),
    .A2(_163_),
    .B1(_169_),
    .Y(_056_));
 sky130_fd_sc_hd__inv_1 _358_ (.A(\gpio[19] ),
    .Y(_170_));
 sky130_fd_sc_hd__o21ai_0 _359_ (.A1(net203),
    .A2(_163_),
    .B1(_074_),
    .Y(_171_));
 sky130_fd_sc_hd__a21oi_1 _360_ (.A1(_170_),
    .A2(_163_),
    .B1(_171_),
    .Y(_057_));
 sky130_fd_sc_hd__inv_1 _361_ (.A(\gpio[20] ),
    .Y(_172_));
 sky130_fd_sc_hd__o21ai_0 _363_ (.A1(net199),
    .A2(_163_),
    .B1(_074_),
    .Y(_174_));
 sky130_fd_sc_hd__a21oi_1 _364_ (.A1(_172_),
    .A2(net942),
    .B1(_174_),
    .Y(_058_));
 sky130_fd_sc_hd__inv_1 _365_ (.A(\gpio[21] ),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _366_ (.A1(net196),
    .A2(_163_),
    .B1(_074_),
    .Y(_176_));
 sky130_fd_sc_hd__a21oi_1 _367_ (.A1(_175_),
    .A2(_163_),
    .B1(_176_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_1 _368_ (.A(\gpio[22] ),
    .Y(_177_));
 sky130_fd_sc_hd__o21ai_0 _369_ (.A1(net192),
    .A2(_163_),
    .B1(_074_),
    .Y(_178_));
 sky130_fd_sc_hd__a21oi_1 _370_ (.A1(_177_),
    .A2(_163_),
    .B1(_178_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_1 _371_ (.A(\gpio[23] ),
    .Y(_179_));
 sky130_fd_sc_hd__o21ai_0 _372_ (.A1(net190),
    .A2(_163_),
    .B1(_074_),
    .Y(_180_));
 sky130_fd_sc_hd__a21oi_1 _373_ (.A1(_179_),
    .A2(net942),
    .B1(_180_),
    .Y(_061_));
 sky130_fd_sc_hd__inv_1 _374_ (.A(\gpio[0] ),
    .Y(_181_));
 sky130_fd_sc_hd__nand4_4 _375_ (.A(net565),
    .B(net718),
    .C(net702),
    .D(_086_),
    .Y(_182_));
 sky130_fd_sc_hd__o21ai_0 _377_ (.A1(net296),
    .A2(_182_),
    .B1(_074_),
    .Y(_184_));
 sky130_fd_sc_hd__a21oi_1 _378_ (.A1(_181_),
    .A2(net703),
    .B1(_184_),
    .Y(_063_));
 sky130_fd_sc_hd__inv_1 _379_ (.A(net4),
    .Y(_185_));
 sky130_fd_sc_hd__o21ai_0 _380_ (.A1(net278),
    .A2(net703),
    .B1(_074_),
    .Y(_186_));
 sky130_fd_sc_hd__a21oi_1 _381_ (.A1(_185_),
    .A2(net703),
    .B1(_186_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_1 _382_ (.A(net5),
    .Y(_187_));
 sky130_fd_sc_hd__o21ai_0 _383_ (.A1(net274),
    .A2(net703),
    .B1(_074_),
    .Y(_188_));
 sky130_fd_sc_hd__a21oi_1 _384_ (.A1(_187_),
    .A2(net703),
    .B1(_188_),
    .Y(_065_));
 sky130_fd_sc_hd__inv_1 _385_ (.A(net6),
    .Y(_189_));
 sky130_fd_sc_hd__o21ai_0 _386_ (.A1(net267),
    .A2(_182_),
    .B1(_074_),
    .Y(_190_));
 sky130_fd_sc_hd__a21oi_1 _387_ (.A1(_189_),
    .A2(_182_),
    .B1(_190_),
    .Y(_066_));
 sky130_fd_sc_hd__inv_1 _388_ (.A(net7),
    .Y(_191_));
 sky130_fd_sc_hd__o21ai_0 _389_ (.A1(net265),
    .A2(_182_),
    .B1(_074_),
    .Y(_192_));
 sky130_fd_sc_hd__a21oi_1 _390_ (.A1(_191_),
    .A2(_182_),
    .B1(_192_),
    .Y(_067_));
 sky130_fd_sc_hd__inv_1 _391_ (.A(net8),
    .Y(_193_));
 sky130_fd_sc_hd__o21ai_0 _392_ (.A1(net263),
    .A2(_182_),
    .B1(_074_),
    .Y(_194_));
 sky130_fd_sc_hd__a21oi_1 _393_ (.A1(_193_),
    .A2(_182_),
    .B1(_194_),
    .Y(_068_));
 sky130_fd_sc_hd__o21ai_0 _394_ (.A1(net256),
    .A2(net703),
    .B1(_074_),
    .Y(_195_));
 sky130_fd_sc_hd__a21oi_1 _395_ (.A1(net10),
    .A2(net703),
    .B1(_195_),
    .Y(_069_));
 sky130_fd_sc_hd__o21ai_0 _396_ (.A1(net253),
    .A2(_182_),
    .B1(_074_),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_1 _397_ (.A1(net9),
    .A2(net703),
    .B1(_196_),
    .Y(_070_));
 sky130_fd_sc_hd__dfxtp_1 _398_ (.CLK(clknet_leaf_62_clk),
    .D(_006_),
    .Q(\gpio[8] ));
 sky130_fd_sc_hd__dfxtp_1 _399_ (.CLK(clknet_leaf_82_clk),
    .D(_007_),
    .Q(\gpio[9] ));
 sky130_fd_sc_hd__dfxtp_1 _400_ (.CLK(clknet_leaf_82_clk),
    .D(_008_),
    .Q(\gpio[10] ));
 sky130_fd_sc_hd__dfxtp_1 _401_ (.CLK(clknet_leaf_83_clk),
    .D(_009_),
    .Q(\gpio[11] ));
 sky130_fd_sc_hd__dfxtp_1 _402_ (.CLK(clknet_leaf_83_clk),
    .D(_010_),
    .Q(\gpio[12] ));
 sky130_fd_sc_hd__dfxtp_1 _403_ (.CLK(clknet_leaf_83_clk),
    .D(_011_),
    .Q(\gpio[13] ));
 sky130_fd_sc_hd__dfxtp_1 _404_ (.CLK(clknet_leaf_82_clk),
    .D(_012_),
    .Q(\gpio[14] ));
 sky130_fd_sc_hd__dfxtp_1 _405_ (.CLK(clknet_leaf_84_clk),
    .D(_013_),
    .Q(\gpio[15] ));
 sky130_fd_sc_hd__dfxtp_1 _406_ (.CLK(clknet_leaf_83_clk),
    .D(_014_),
    .Q(\iomem_rdata[0] ));
 sky130_fd_sc_hd__dfxtp_1 _407_ (.CLK(clknet_leaf_82_clk),
    .D(net770),
    .Q(\iomem_rdata[1] ));
 sky130_fd_sc_hd__dfxtp_1 _408_ (.CLK(clknet_leaf_82_clk),
    .D(net759),
    .Q(\iomem_rdata[2] ));
 sky130_fd_sc_hd__dfxtp_1 _409_ (.CLK(clknet_leaf_83_clk),
    .D(_017_),
    .Q(\iomem_rdata[3] ));
 sky130_fd_sc_hd__dfxtp_1 _410_ (.CLK(clknet_leaf_83_clk),
    .D(_018_),
    .Q(\iomem_rdata[4] ));
 sky130_fd_sc_hd__dfxtp_1 _411_ (.CLK(clknet_leaf_83_clk),
    .D(_019_),
    .Q(\iomem_rdata[5] ));
 sky130_fd_sc_hd__dfxtp_1 _412_ (.CLK(clknet_leaf_74_clk),
    .D(_020_),
    .Q(\iomem_rdata[6] ));
 sky130_fd_sc_hd__dfxtp_1 _413_ (.CLK(clknet_leaf_62_clk),
    .D(_021_),
    .Q(\iomem_rdata[7] ));
 sky130_fd_sc_hd__dfxtp_1 _414_ (.CLK(clknet_leaf_62_clk),
    .D(_022_),
    .Q(\iomem_rdata[8] ));
 sky130_fd_sc_hd__dfxtp_1 _415_ (.CLK(clknet_leaf_82_clk),
    .D(_023_),
    .Q(\iomem_rdata[9] ));
 sky130_fd_sc_hd__dfxtp_1 _416_ (.CLK(clknet_leaf_83_clk),
    .D(_024_),
    .Q(\iomem_rdata[10] ));
 sky130_fd_sc_hd__dfxtp_1 _417_ (.CLK(clknet_leaf_83_clk),
    .D(_025_),
    .Q(\iomem_rdata[11] ));
 sky130_fd_sc_hd__dfxtp_1 _418_ (.CLK(clknet_leaf_84_clk),
    .D(_026_),
    .Q(\iomem_rdata[12] ));
 sky130_fd_sc_hd__dfxtp_1 _419_ (.CLK(clknet_leaf_83_clk),
    .D(_027_),
    .Q(\iomem_rdata[13] ));
 sky130_fd_sc_hd__dfxtp_1 _420_ (.CLK(clknet_leaf_82_clk),
    .D(_028_),
    .Q(\iomem_rdata[14] ));
 sky130_fd_sc_hd__dfxtp_1 _421_ (.CLK(clknet_leaf_84_clk),
    .D(_029_),
    .Q(\iomem_rdata[15] ));
 sky130_fd_sc_hd__dfxtp_1 _422_ (.CLK(clknet_leaf_84_clk),
    .D(_030_),
    .Q(\iomem_rdata[16] ));
 sky130_fd_sc_hd__dfxtp_1 _423_ (.CLK(clknet_leaf_80_clk),
    .D(_031_),
    .Q(\iomem_rdata[17] ));
 sky130_fd_sc_hd__dfxtp_1 _424_ (.CLK(clknet_leaf_80_clk),
    .D(_032_),
    .Q(\iomem_rdata[18] ));
 sky130_fd_sc_hd__dfxtp_1 _425_ (.CLK(clknet_leaf_85_clk),
    .D(_033_),
    .Q(\iomem_rdata[19] ));
 sky130_fd_sc_hd__dfxtp_1 _426_ (.CLK(clknet_leaf_84_clk),
    .D(_034_),
    .Q(\iomem_rdata[20] ));
 sky130_fd_sc_hd__dfxtp_1 _427_ (.CLK(clknet_leaf_85_clk),
    .D(_035_),
    .Q(\iomem_rdata[21] ));
 sky130_fd_sc_hd__dfxtp_1 _428_ (.CLK(clknet_leaf_80_clk),
    .D(_036_),
    .Q(\iomem_rdata[22] ));
 sky130_fd_sc_hd__dfxtp_1 _429_ (.CLK(clknet_leaf_84_clk),
    .D(_037_),
    .Q(\iomem_rdata[23] ));
 sky130_fd_sc_hd__dfxtp_1 _430_ (.CLK(clknet_leaf_80_clk),
    .D(_038_),
    .Q(\iomem_rdata[24] ));
 sky130_fd_sc_hd__dfxtp_1 _431_ (.CLK(clknet_leaf_85_clk),
    .D(_039_),
    .Q(\iomem_rdata[25] ));
 sky130_fd_sc_hd__dfxtp_1 _432_ (.CLK(clknet_leaf_80_clk),
    .D(_040_),
    .Q(\iomem_rdata[26] ));
 sky130_fd_sc_hd__dfxtp_1 _433_ (.CLK(clknet_leaf_89_clk),
    .D(_041_),
    .Q(\iomem_rdata[27] ));
 sky130_fd_sc_hd__dfxtp_1 _434_ (.CLK(clknet_leaf_85_clk),
    .D(_042_),
    .Q(\iomem_rdata[28] ));
 sky130_fd_sc_hd__dfxtp_1 _435_ (.CLK(clknet_leaf_85_clk),
    .D(_043_),
    .Q(\iomem_rdata[29] ));
 sky130_fd_sc_hd__dfxtp_1 _436_ (.CLK(clknet_leaf_81_clk),
    .D(net706),
    .Q(\iomem_rdata[30] ));
 sky130_fd_sc_hd__dfxtp_1 _437_ (.CLK(clknet_leaf_85_clk),
    .D(_045_),
    .Q(\iomem_rdata[31] ));
 sky130_fd_sc_hd__dfxtp_1 _438_ (.CLK(clknet_leaf_91_clk),
    .D(_046_),
    .Q(\gpio[24] ));
 sky130_fd_sc_hd__dfxtp_1 _439_ (.CLK(clknet_leaf_85_clk),
    .D(_047_),
    .Q(\gpio[25] ));
 sky130_fd_sc_hd__dfxtp_1 _440_ (.CLK(clknet_leaf_80_clk),
    .D(_048_),
    .Q(\gpio[26] ));
 sky130_fd_sc_hd__dfxtp_1 _441_ (.CLK(clknet_leaf_89_clk),
    .D(_049_),
    .Q(\gpio[27] ));
 sky130_fd_sc_hd__dfxtp_1 _442_ (.CLK(clknet_leaf_91_clk),
    .D(_050_),
    .Q(\gpio[28] ));
 sky130_fd_sc_hd__dfxtp_1 _443_ (.CLK(clknet_leaf_85_clk),
    .D(_051_),
    .Q(\gpio[29] ));
 sky130_fd_sc_hd__dfxtp_2 _444_ (.CLK(clknet_leaf_85_clk),
    .D(_052_),
    .Q(\gpio[30] ));
 sky130_fd_sc_hd__dfxtp_1 _445_ (.CLK(clknet_leaf_89_clk),
    .D(_053_),
    .Q(\gpio[31] ));
 sky130_fd_sc_hd__dfxtp_1 _446_ (.CLK(clknet_leaf_84_clk),
    .D(_054_),
    .Q(\gpio[16] ));
 sky130_fd_sc_hd__dfxtp_1 _447_ (.CLK(clknet_leaf_80_clk),
    .D(_055_),
    .Q(\gpio[17] ));
 sky130_fd_sc_hd__dfxtp_1 _448_ (.CLK(clknet_leaf_80_clk),
    .D(_056_),
    .Q(\gpio[18] ));
 sky130_fd_sc_hd__dfxtp_1 _449_ (.CLK(clknet_leaf_85_clk),
    .D(_057_),
    .Q(\gpio[19] ));
 sky130_fd_sc_hd__dfxtp_1 _450_ (.CLK(clknet_leaf_84_clk),
    .D(_058_),
    .Q(\gpio[20] ));
 sky130_fd_sc_hd__dfxtp_1 _451_ (.CLK(clknet_leaf_85_clk),
    .D(_059_),
    .Q(\gpio[21] ));
 sky130_fd_sc_hd__dfxtp_1 _452_ (.CLK(clknet_leaf_80_clk),
    .D(_060_),
    .Q(\gpio[22] ));
 sky130_fd_sc_hd__dfxtp_1 _453_ (.CLK(clknet_leaf_84_clk),
    .D(_061_),
    .Q(\gpio[23] ));
 sky130_fd_sc_hd__dfxtp_1 _454_ (.CLK(clknet_leaf_85_clk),
    .D(_062_),
    .Q(iomem_ready));
 sky130_fd_sc_hd__dfxtp_1 _455_ (.CLK(clknet_leaf_61_clk),
    .D(_063_),
    .Q(\gpio[0] ));
 sky130_fd_sc_hd__dfxtp_4 _456_ (.CLK(clknet_leaf_81_clk),
    .D(_064_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_4 _457_ (.CLK(clknet_leaf_82_clk),
    .D(_065_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_4 _458_ (.CLK(clknet_leaf_83_clk),
    .D(_066_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_4 _459_ (.CLK(clknet_leaf_83_clk),
    .D(_067_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_4 _460_ (.CLK(clknet_leaf_83_clk),
    .D(_068_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _461_ (.CLK(clknet_leaf_74_clk),
    .D(_069_),
    .Q(\gpio[6] ));
 sky130_fd_sc_hd__dfxtp_1 _462_ (.CLK(clknet_leaf_61_clk),
    .D(_070_),
    .Q(\gpio[7] ));
 sky130_fd_sc_hd__dfxtp_1 _463_ (.CLK(clknet_leaf_62_clk),
    .D(_000_),
    .Q(\reset_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _464_ (.CLK(clknet_leaf_62_clk),
    .D(_001_),
    .Q(\reset_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _465_ (.CLK(clknet_leaf_62_clk),
    .D(_002_),
    .Q(\reset_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _466_ (.CLK(clknet_leaf_62_clk),
    .D(_003_),
    .Q(\reset_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _467_ (.CLK(clknet_leaf_82_clk),
    .D(_004_),
    .Q(\reset_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _468_ (.CLK(clknet_leaf_62_clk),
    .D(_005_),
    .Q(\reset_cnt[5] ));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06653__419  (.LO(net419));
 sky130_fd_sc_hd__nor4_1 \soc/_233_  (.A(\iomem_addr[22] ),
    .B(\iomem_addr[19] ),
    .C(net724),
    .D(net779),
    .Y(\soc/_013_ ));
 sky130_fd_sc_hd__nor4_1 \soc/_234_  (.A(\iomem_addr[24] ),
    .B(\iomem_addr[21] ),
    .C(\iomem_addr[20] ),
    .D(net694),
    .Y(\soc/_014_ ));
 sky130_fd_sc_hd__nor4_1 \soc/_235_  (.A(\iomem_addr[13] ),
    .B(net771),
    .C(net713),
    .D(net708),
    .Y(\soc/_015_ ));
 sky130_fd_sc_hd__nor3_1 \soc/_236_  (.A(net736),
    .B(net744),
    .C(net714),
    .Y(\soc/_016_ ));
 sky130_fd_sc_hd__nand4_4 \soc/_237_  (.A(net725),
    .B(\soc/_014_ ),
    .C(\soc/_015_ ),
    .D(\soc/_016_ ),
    .Y(\soc/_017_ ));
 sky130_fd_sc_hd__nor2_2 \soc/_238_  (.A(net717),
    .B(net739),
    .Y(\soc/_018_ ));
 sky130_fd_sc_hd__nor4_4 \soc/_239_  (.A(\iomem_addr[28] ),
    .B(net701),
    .C(net809),
    .D(net763),
    .Y(\soc/_019_ ));
 sky130_fd_sc_hd__nor2_1 \soc/_240_  (.A(net521),
    .B(net515),
    .Y(\soc/_020_ ));
 sky130_fd_sc_hd__nand4_4 \soc/_241_  (.A(net492),
    .B(net740),
    .C(net764),
    .D(\soc/_020_ ),
    .Y(\soc/_021_ ));
 sky130_fd_sc_hd__nor4_1 \soc/_242_  (.A(net497),
    .B(net367),
    .C(net501),
    .D(net378),
    .Y(\soc/_022_ ));
 sky130_fd_sc_hd__nor4b_1 \soc/_243_  (.A(net448),
    .B(net449),
    .C(net391),
    .D_N(net386),
    .Y(\soc/_023_ ));
 sky130_fd_sc_hd__nand3_1 \soc/_244_  (.A(net903),
    .B(\soc/_022_ ),
    .C(\soc/_023_ ),
    .Y(\soc/_024_ ));
 sky130_fd_sc_hd__nor3_4 \soc/_245_  (.A(net726),
    .B(net741),
    .C(\soc/_024_ ),
    .Y(\soc/_025_ ));
 sky130_fd_sc_hd__inv_1 \soc/_246_  (.A(net138),
    .Y(\soc/_026_ ));
 sky130_fd_sc_hd__inv_1 \soc/_247_  (.A(net492),
    .Y(\soc/_027_ ));
 sky130_fd_sc_hd__inv_1 \soc/_248_  (.A(net808),
    .Y(\soc/_028_ ));
 sky130_fd_sc_hd__inv_1 \soc/_249_  (.A(net903),
    .Y(\soc/_029_ ));
 sky130_fd_sc_hd__a311oi_4 \soc/_250_  (.A1(\soc/_027_ ),
    .A2(net740),
    .A3(net764),
    .B1(\soc/_028_ ),
    .C1(\soc/_029_ ),
    .Y(\soc/_030_ ));
 sky130_fd_sc_hd__or3_1 \soc/_251_  (.A(net109),
    .B(\soc/ram_ready ),
    .C(net146),
    .X(\soc/_031_ ));
 sky130_fd_sc_hd__nor3_1 \soc/_252_  (.A(net450),
    .B(net451),
    .C(net385),
    .Y(\soc/_032_ ));
 sky130_fd_sc_hd__nand4_2 \soc/_253_  (.A(net903),
    .B(net391),
    .C(\soc/_022_ ),
    .D(\soc/_032_ ),
    .Y(\soc/_033_ ));
 sky130_fd_sc_hd__nor3_4 \soc/_254_  (.A(net726),
    .B(net741),
    .C(net904),
    .Y(\soc/_034_ ));
 sky130_fd_sc_hd__nand4b_1 \soc/_256_  (.A_N(net391),
    .B(\soc/_022_ ),
    .C(\soc/_032_ ),
    .D(net903),
    .Y(\soc/_036_ ));
 sky130_fd_sc_hd__nor3_1 \soc/_257_  (.A(net726),
    .B(net741),
    .C(\soc/_036_ ),
    .Y(\soc/_037_ ));
 sky130_fd_sc_hd__nor3_2 \soc/_259_  (.A(\soc/_031_ ),
    .B(net906),
    .C(net743),
    .Y(\soc/_039_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_260_  (.A1(\soc/simpleuart_reg_dat_wait ),
    .A2(\soc/_026_ ),
    .B1(net907),
    .Y(\soc/mem_ready ));
 sky130_fd_sc_hd__nand2_1 \soc/_261_  (.A(net740),
    .B(net764),
    .Y(\soc/_040_ ));
 sky130_fd_sc_hd__or4_4 \soc/_262_  (.A(\soc/_029_ ),
    .B(net492),
    .C(net765),
    .D(net726),
    .X(\soc/_041_ ));
 sky130_fd_sc_hd__nor2_1 \soc/_263_  (.A(\soc/mem_ready ),
    .B(net493),
    .Y(\soc/_000_ ));
 sky130_fd_sc_hd__nor4_2 \soc/_264_  (.A(net563),
    .B(net568),
    .C(net545),
    .D(net577),
    .Y(\soc/_042_ ));
 sky130_fd_sc_hd__nor3_2 \soc/_265_  (.A(net908),
    .B(net767),
    .C(\soc/_042_ ),
    .Y(\soc/_003_ ));
 sky130_fd_sc_hd__and2_0 \soc/_267_  (.A(net138),
    .B(\soc/_042_ ),
    .X(\soc/_002_ ));
 sky130_fd_sc_hd__nor2_1 \soc/_268_  (.A(net492),
    .B(\soc/_040_ ),
    .Y(\soc/_044_ ));
 sky130_fd_sc_hd__and3_2 \soc/_269_  (.A(\soc/mem_valid ),
    .B(\soc/_044_ ),
    .C(net726),
    .X(\soc/_001_ ));
 sky130_fd_sc_hd__nor2_1 \soc/_270_  (.A(\soc/_029_ ),
    .B(\soc/_044_ ),
    .Y(iomem_valid));
 sky130_fd_sc_hd__and2_2 \soc/_271_  (.A(net410),
    .B(net136),
    .X(\soc/_008_ ));
 sky130_fd_sc_hd__and2_1 \soc/_272_  (.A(net406),
    .B(net136),
    .X(\soc/_009_ ));
 sky130_fd_sc_hd__and2_2 \soc/_273_  (.A(net402),
    .B(net136),
    .X(\soc/_010_ ));
 sky130_fd_sc_hd__and2_2 \soc/_274_  (.A(net545),
    .B(net136),
    .X(\soc/_011_ ));
 sky130_fd_sc_hd__and2_4 \soc/_275_  (.A(net411),
    .B(net135),
    .X(\soc/_004_ ));
 sky130_fd_sc_hd__and2_2 \soc/_276_  (.A(net406),
    .B(net135),
    .X(\soc/_005_ ));
 sky130_fd_sc_hd__and2_2 \soc/_277_  (.A(net402),
    .B(net135),
    .X(\soc/_006_ ));
 sky130_fd_sc_hd__and2_0 \soc/_278_  (.A(net400),
    .B(net135),
    .X(\soc/_007_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/_283_  (.A1(\soc/simpleuart_reg_div_do[0] ),
    .A2(net136),
    .B1(net134),
    .B2(flash_io0),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[0] ),
    .Y(\soc/_049_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_287_  (.A1(net415),
    .A2(\soc/ram_rdata[0] ),
    .B1(net108),
    .Y(\soc/_053_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_288_  (.A1(net415),
    .A2(\soc/_049_ ),
    .B1(\soc/_053_ ),
    .Y(\soc/_054_ ));
 sky130_fd_sc_hd__inv_1 \soc/_290_  (.A(\soc/spimem_rdata[0] ),
    .Y(\soc/_056_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_292_  (.A1(net111),
    .A2(\soc/_056_ ),
    .B1(net149),
    .Y(\soc/_058_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_293_  (.A1(\iomem_rdata[0] ),
    .A2(net149),
    .B1(\soc/_054_ ),
    .B2(\soc/_058_ ),
    .X(\soc/mem_rdata[0] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_294_  (.A1(\soc/simpleuart_reg_div_do[1] ),
    .A2(net136),
    .B1(net134),
    .B2(flash_io1),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[1] ),
    .Y(\soc/_059_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_295_  (.A1(net415),
    .A2(\soc/ram_rdata[1] ),
    .B1(net108),
    .Y(\soc/_060_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_296_  (.A1(net415),
    .A2(\soc/_059_ ),
    .B1(\soc/_060_ ),
    .Y(\soc/_061_ ));
 sky130_fd_sc_hd__inv_1 \soc/_297_  (.A(\soc/spimem_rdata[1] ),
    .Y(\soc/_062_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_298_  (.A1(net111),
    .A2(\soc/_062_ ),
    .B1(net146),
    .Y(\soc/_063_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_299_  (.A1(\iomem_rdata[1] ),
    .A2(net146),
    .B1(\soc/_061_ ),
    .B2(\soc/_063_ ),
    .X(\soc/mem_rdata[1] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_300_  (.A1(\soc/simpleuart_reg_div_do[2] ),
    .A2(net136),
    .B1(net134),
    .B2(flash_io2),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[2] ),
    .Y(\soc/_064_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_301_  (.A1(net415),
    .A2(\soc/ram_rdata[2] ),
    .B1(net108),
    .Y(\soc/_065_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_302_  (.A1(net415),
    .A2(\soc/_064_ ),
    .B1(\soc/_065_ ),
    .Y(\soc/_066_ ));
 sky130_fd_sc_hd__inv_1 \soc/_303_  (.A(\soc/spimem_rdata[2] ),
    .Y(\soc/_067_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_304_  (.A1(net111),
    .A2(\soc/_067_ ),
    .B1(net147),
    .Y(\soc/_068_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_305_  (.A1(\iomem_rdata[2] ),
    .A2(net147),
    .B1(\soc/_066_ ),
    .B2(\soc/_068_ ),
    .X(\soc/mem_rdata[2] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_306_  (.A1(\soc/simpleuart_reg_div_do[3] ),
    .A2(net136),
    .B1(net134),
    .B2(flash_io3),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[3] ),
    .Y(\soc/_069_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_307_  (.A1(net415),
    .A2(\soc/ram_rdata[3] ),
    .B1(net108),
    .Y(\soc/_070_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_308_  (.A1(net415),
    .A2(\soc/_069_ ),
    .B1(\soc/_070_ ),
    .Y(\soc/_071_ ));
 sky130_fd_sc_hd__inv_1 \soc/_309_  (.A(\soc/spimem_rdata[3] ),
    .Y(\soc/_072_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_310_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_072_ ),
    .B1(net147),
    .Y(\soc/_073_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_311_  (.A1(\iomem_rdata[3] ),
    .A2(net147),
    .B1(\soc/_071_ ),
    .B2(\soc/_073_ ),
    .X(\soc/mem_rdata[3] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_312_  (.A1(\soc/simpleuart_reg_div_do[4] ),
    .A2(net136),
    .B1(net134),
    .B2(net2),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[4] ),
    .Y(\soc/_074_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_313_  (.A1(net415),
    .A2(\soc/ram_rdata[4] ),
    .B1(net108),
    .Y(\soc/_075_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_314_  (.A1(net415),
    .A2(\soc/_074_ ),
    .B1(\soc/_075_ ),
    .Y(\soc/_076_ ));
 sky130_fd_sc_hd__inv_1 \soc/_315_  (.A(\soc/spimem_rdata[4] ),
    .Y(\soc/_077_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_316_  (.A1(net110),
    .A2(\soc/_077_ ),
    .B1(net149),
    .Y(\soc/_078_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_317_  (.A1(\iomem_rdata[4] ),
    .A2(net149),
    .B1(\soc/_076_ ),
    .B2(\soc/_078_ ),
    .X(\soc/mem_rdata[4] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_320_  (.A1(\soc/simpleuart_reg_div_do[5] ),
    .A2(net136),
    .B1(net134),
    .B2(net3),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[5] ),
    .Y(\soc/_081_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_321_  (.A1(net415),
    .A2(\soc/ram_rdata[5] ),
    .B1(net108),
    .Y(\soc/_082_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_322_  (.A1(net415),
    .A2(\soc/_081_ ),
    .B1(\soc/_082_ ),
    .Y(\soc/_083_ ));
 sky130_fd_sc_hd__inv_1 \soc/_323_  (.A(\soc/spimem_rdata[5] ),
    .Y(\soc/_084_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_324_  (.A1(net110),
    .A2(\soc/_084_ ),
    .B1(net149),
    .Y(\soc/_085_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_325_  (.A1(\iomem_rdata[5] ),
    .A2(net149),
    .B1(\soc/_083_ ),
    .B2(\soc/_085_ ),
    .X(\soc/mem_rdata[5] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_326_  (.A1(\soc/simpleuart_reg_div_do[6] ),
    .A2(net136),
    .B1(net134),
    .B2(net458),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[6] ),
    .Y(\soc/_086_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_327_  (.A1(net415),
    .A2(\soc/ram_rdata[6] ),
    .B1(net108),
    .Y(\soc/_087_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_328_  (.A1(net415),
    .A2(\soc/_086_ ),
    .B1(\soc/_087_ ),
    .Y(\soc/_088_ ));
 sky130_fd_sc_hd__inv_1 \soc/_329_  (.A(\soc/spimem_rdata[6] ),
    .Y(\soc/_089_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_330_  (.A1(net111),
    .A2(\soc/_089_ ),
    .B1(net146),
    .Y(\soc/_090_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_331_  (.A1(\iomem_rdata[6] ),
    .A2(net146),
    .B1(\soc/_088_ ),
    .B2(\soc/_090_ ),
    .X(\soc/mem_rdata[6] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_332_  (.A1(\soc/simpleuart_reg_div_do[7] ),
    .A2(net136),
    .B1(net134),
    .B2(net459),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[7] ),
    .Y(\soc/_091_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_333_  (.A1(net415),
    .A2(\soc/ram_rdata[7] ),
    .B1(net108),
    .Y(\soc/_092_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_334_  (.A1(net415),
    .A2(\soc/_091_ ),
    .B1(\soc/_092_ ),
    .Y(\soc/_093_ ));
 sky130_fd_sc_hd__inv_1 \soc/_335_  (.A(\soc/spimem_rdata[7] ),
    .Y(\soc/_094_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_336_  (.A1(net111),
    .A2(\soc/_094_ ),
    .B1(net149),
    .Y(\soc/_095_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_337_  (.A1(\iomem_rdata[7] ),
    .A2(net149),
    .B1(\soc/_093_ ),
    .B2(\soc/_095_ ),
    .X(\soc/mem_rdata[7] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_339_  (.A1(\soc/simpleuart_reg_div_do[8] ),
    .A2(net137),
    .B1(net134),
    .B2(flash_io0_oe),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_097_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_342_  (.A1(net415),
    .A2(\soc/ram_rdata[8] ),
    .B1(net109),
    .Y(\soc/_100_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_343_  (.A1(net415),
    .A2(\soc/_097_ ),
    .B1(\soc/_100_ ),
    .Y(\soc/_101_ ));
 sky130_fd_sc_hd__inv_1 \soc/_344_  (.A(\soc/spimem_rdata[8] ),
    .Y(\soc/_102_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_346_  (.A1(net111),
    .A2(\soc/_102_ ),
    .B1(net149),
    .Y(\soc/_104_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_347_  (.A1(\iomem_rdata[8] ),
    .A2(net149),
    .B1(\soc/_101_ ),
    .B2(\soc/_104_ ),
    .X(\soc/mem_rdata[8] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_348_  (.A1(\soc/simpleuart_reg_div_do[9] ),
    .A2(net137),
    .B1(net134),
    .B2(flash_io1_oe),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_105_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_349_  (.A1(net415),
    .A2(\soc/ram_rdata[9] ),
    .B1(net109),
    .Y(\soc/_106_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_350_  (.A1(net415),
    .A2(\soc/_105_ ),
    .B1(\soc/_106_ ),
    .Y(\soc/_107_ ));
 sky130_fd_sc_hd__inv_1 \soc/_351_  (.A(\soc/spimem_rdata[9] ),
    .Y(\soc/_108_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_352_  (.A1(net111),
    .A2(\soc/_108_ ),
    .B1(net147),
    .Y(\soc/_109_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_353_  (.A1(\iomem_rdata[9] ),
    .A2(net147),
    .B1(\soc/_107_ ),
    .B2(\soc/_109_ ),
    .X(\soc/mem_rdata[9] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_356_  (.A1(\soc/simpleuart_reg_div_do[10] ),
    .A2(net137),
    .B1(net134),
    .B2(flash_io2_oe),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_112_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_357_  (.A1(net415),
    .A2(\soc/ram_rdata[10] ),
    .B1(net109),
    .Y(\soc/_113_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_358_  (.A1(net415),
    .A2(\soc/_112_ ),
    .B1(\soc/_113_ ),
    .Y(\soc/_114_ ));
 sky130_fd_sc_hd__inv_1 \soc/_360_  (.A(\soc/spimem_rdata[10] ),
    .Y(\soc/_116_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_361_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_116_ ),
    .B1(net147),
    .Y(\soc/_117_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_362_  (.A1(\iomem_rdata[10] ),
    .A2(net147),
    .B1(\soc/_114_ ),
    .B2(\soc/_117_ ),
    .X(\soc/mem_rdata[10] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_363_  (.A1(\soc/simpleuart_reg_div_do[11] ),
    .A2(net137),
    .B1(net134),
    .B2(flash_io3_oe),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_118_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_364_  (.A1(net415),
    .A2(\soc/ram_rdata[11] ),
    .B1(net109),
    .Y(\soc/_119_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_365_  (.A1(net415),
    .A2(\soc/_118_ ),
    .B1(\soc/_119_ ),
    .Y(\soc/_120_ ));
 sky130_fd_sc_hd__inv_1 \soc/_366_  (.A(\soc/spimem_rdata[11] ),
    .Y(\soc/_121_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_367_  (.A1(net110),
    .A2(\soc/_121_ ),
    .B1(net149),
    .Y(\soc/_122_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_368_  (.A1(\iomem_rdata[11] ),
    .A2(net149),
    .B1(\soc/_120_ ),
    .B2(\soc/_122_ ),
    .X(\soc/mem_rdata[11] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_369_  (.A1(\soc/simpleuart_reg_div_do[12] ),
    .A2(net137),
    .B1(net134),
    .B2(net460),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_123_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/_370_  (.A1(net415),
    .A2(\soc/ram_rdata[12] ),
    .B1(net108),
    .Y(\soc/_124_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_371_  (.A1(net415),
    .A2(\soc/_123_ ),
    .B1(\soc/_124_ ),
    .Y(\soc/_125_ ));
 sky130_fd_sc_hd__inv_1 \soc/_372_  (.A(\soc/spimem_rdata[12] ),
    .Y(\soc/_126_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_373_  (.A1(net110),
    .A2(\soc/_126_ ),
    .B1(net149),
    .Y(\soc/_127_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_374_  (.A1(\iomem_rdata[12] ),
    .A2(\soc/_030_ ),
    .B1(\soc/_125_ ),
    .B2(\soc/_127_ ),
    .X(\soc/mem_rdata[12] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_375_  (.A1(\soc/simpleuart_reg_div_do[13] ),
    .A2(net137),
    .B1(net134),
    .B2(net461),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_128_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_376_  (.A1(net415),
    .A2(\soc/ram_rdata[13] ),
    .B1(net109),
    .Y(\soc/_129_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_377_  (.A1(net415),
    .A2(\soc/_128_ ),
    .B1(\soc/_129_ ),
    .Y(\soc/_130_ ));
 sky130_fd_sc_hd__inv_1 \soc/_378_  (.A(\soc/spimem_rdata[13] ),
    .Y(\soc/_131_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_379_  (.A1(net110),
    .A2(\soc/_131_ ),
    .B1(net149),
    .Y(\soc/_132_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_380_  (.A1(\iomem_rdata[13] ),
    .A2(net149),
    .B1(\soc/_130_ ),
    .B2(\soc/_132_ ),
    .X(\soc/mem_rdata[13] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_381_  (.A1(\soc/simpleuart_reg_div_do[14] ),
    .A2(net136),
    .B1(net134),
    .B2(net462),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_133_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_382_  (.A1(net415),
    .A2(\soc/ram_rdata[14] ),
    .B1(net108),
    .Y(\soc/_134_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_383_  (.A1(net415),
    .A2(\soc/_133_ ),
    .B1(\soc/_134_ ),
    .Y(\soc/_135_ ));
 sky130_fd_sc_hd__inv_1 \soc/_384_  (.A(\soc/spimem_rdata[14] ),
    .Y(\soc/_136_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_385_  (.A1(net111),
    .A2(\soc/_136_ ),
    .B1(net146),
    .Y(\soc/_137_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_386_  (.A1(\iomem_rdata[14] ),
    .A2(net146),
    .B1(\soc/_135_ ),
    .B2(\soc/_137_ ),
    .X(\soc/mem_rdata[14] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_389_  (.A1(\soc/simpleuart_reg_div_do[15] ),
    .A2(net136),
    .B1(net134),
    .B2(net463),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_140_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_390_  (.A1(net415),
    .A2(\soc/ram_rdata[15] ),
    .B1(net108),
    .Y(\soc/_141_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_391_  (.A1(net415),
    .A2(\soc/_140_ ),
    .B1(\soc/_141_ ),
    .Y(\soc/_142_ ));
 sky130_fd_sc_hd__inv_1 \soc/_392_  (.A(\soc/spimem_rdata[15] ),
    .Y(\soc/_143_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_393_  (.A1(net110),
    .A2(\soc/_143_ ),
    .B1(net149),
    .Y(\soc/_144_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_394_  (.A1(\iomem_rdata[15] ),
    .A2(net149),
    .B1(\soc/_142_ ),
    .B2(\soc/_144_ ),
    .X(\soc/mem_rdata[15] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_395_  (.A1(\soc/simpleuart_reg_div_do[16] ),
    .A2(net137),
    .B1(net135),
    .B2(\soc/spimemio_cfgreg_do[16] ),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_145_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_396_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[16] ),
    .B1(net109),
    .Y(\soc/_146_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_397_  (.A1(\soc/ram_ready ),
    .A2(\soc/_145_ ),
    .B1(\soc/_146_ ),
    .Y(\soc/_147_ ));
 sky130_fd_sc_hd__inv_1 \soc/_398_  (.A(\soc/spimem_rdata[16] ),
    .Y(\soc/_148_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_399_  (.A1(net110),
    .A2(\soc/_148_ ),
    .B1(\soc/_030_ ),
    .Y(\soc/_149_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_400_  (.A1(\iomem_rdata[16] ),
    .A2(\soc/_030_ ),
    .B1(\soc/_147_ ),
    .B2(\soc/_149_ ),
    .X(\soc/mem_rdata[16] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_401_  (.A1(\soc/simpleuart_reg_div_do[17] ),
    .A2(net137),
    .B1(net135),
    .B2(\soc/spimemio_cfgreg_do[17] ),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_150_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_402_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[17] ),
    .B1(net109),
    .Y(\soc/_151_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_403_  (.A1(\soc/ram_ready ),
    .A2(\soc/_150_ ),
    .B1(\soc/_151_ ),
    .Y(\soc/_152_ ));
 sky130_fd_sc_hd__inv_1 \soc/_404_  (.A(\soc/spimem_rdata[17] ),
    .Y(\soc/_153_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_405_  (.A1(net111),
    .A2(\soc/_153_ ),
    .B1(net146),
    .Y(\soc/_154_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_406_  (.A1(net858),
    .A2(net147),
    .B1(\soc/_152_ ),
    .B2(\soc/_154_ ),
    .X(\soc/mem_rdata[17] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_408_  (.A1(\soc/simpleuart_reg_div_do[18] ),
    .A2(net137),
    .B1(net135),
    .B2(\soc/spimemio_cfgreg_do[18] ),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_156_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_411_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[18] ),
    .B1(net109),
    .Y(\soc/_159_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_412_  (.A1(\soc/ram_ready ),
    .A2(\soc/_156_ ),
    .B1(\soc/_159_ ),
    .Y(\soc/_160_ ));
 sky130_fd_sc_hd__inv_1 \soc/_413_  (.A(\soc/spimem_rdata[18] ),
    .Y(\soc/_161_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_415_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_161_ ),
    .B1(net148),
    .Y(\soc/_163_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_416_  (.A1(\iomem_rdata[18] ),
    .A2(net148),
    .B1(\soc/_160_ ),
    .B2(\soc/_163_ ),
    .X(\soc/mem_rdata[18] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_417_  (.A1(\soc/simpleuart_reg_div_do[19] ),
    .A2(\soc/_034_ ),
    .B1(\soc/_037_ ),
    .B2(\soc/spimemio_cfgreg_do[19] ),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_164_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_418_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[19] ),
    .B1(net112),
    .Y(\soc/_165_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_419_  (.A1(\soc/ram_ready ),
    .A2(\soc/_164_ ),
    .B1(\soc/_165_ ),
    .Y(\soc/_166_ ));
 sky130_fd_sc_hd__inv_1 \soc/_420_  (.A(\soc/spimem_rdata[19] ),
    .Y(\soc/_167_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_421_  (.A1(net110),
    .A2(\soc/_167_ ),
    .B1(net150),
    .Y(\soc/_168_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_422_  (.A1(net958),
    .A2(net150),
    .B1(\soc/_166_ ),
    .B2(\soc/_168_ ),
    .X(\soc/mem_rdata[19] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_425_  (.A1(\soc/simpleuart_reg_div_do[20] ),
    .A2(net137),
    .B1(net135),
    .B2(\soc/spimemio/config_cont ),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_171_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_426_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[20] ),
    .B1(net109),
    .Y(\soc/_172_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_427_  (.A1(\soc/ram_ready ),
    .A2(\soc/_171_ ),
    .B1(\soc/_172_ ),
    .Y(\soc/_173_ ));
 sky130_fd_sc_hd__inv_1 \soc/_429_  (.A(\soc/spimem_rdata[20] ),
    .Y(\soc/_175_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_430_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_175_ ),
    .B1(net147),
    .Y(\soc/_176_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_431_  (.A1(\iomem_rdata[20] ),
    .A2(net147),
    .B1(\soc/_173_ ),
    .B2(\soc/_176_ ),
    .X(\soc/mem_rdata[20] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_432_  (.A1(\soc/simpleuart_reg_div_do[21] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(\soc/spimemio/config_qspi ),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_177_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_433_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[21] ),
    .B1(net112),
    .Y(\soc/_178_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_434_  (.A1(\soc/ram_ready ),
    .A2(\soc/_177_ ),
    .B1(\soc/_178_ ),
    .Y(\soc/_179_ ));
 sky130_fd_sc_hd__inv_1 \soc/_435_  (.A(\soc/spimem_rdata[21] ),
    .Y(\soc/_180_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_436_  (.A1(net110),
    .A2(\soc/_180_ ),
    .B1(net150),
    .Y(\soc/_181_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_437_  (.A1(net805),
    .A2(\soc/_030_ ),
    .B1(\soc/_179_ ),
    .B2(\soc/_181_ ),
    .X(\soc/mem_rdata[21] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_438_  (.A1(\soc/simpleuart_reg_div_do[22] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(\soc/spimemio/config_ddr ),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_182_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_439_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[22] ),
    .B1(net112),
    .Y(\soc/_183_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_440_  (.A1(\soc/ram_ready ),
    .A2(\soc/_182_ ),
    .B1(\soc/_183_ ),
    .Y(\soc/_184_ ));
 sky130_fd_sc_hd__inv_1 \soc/_441_  (.A(\soc/spimem_rdata[22] ),
    .Y(\soc/_185_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_442_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_185_ ),
    .B1(net148),
    .Y(\soc/_186_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_443_  (.A1(net859),
    .A2(net148),
    .B1(\soc/_184_ ),
    .B2(\soc/_186_ ),
    .X(\soc/mem_rdata[22] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_444_  (.A1(\soc/simpleuart_reg_div_do[23] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net464),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_187_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_445_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[23] ),
    .B1(net112),
    .Y(\soc/_188_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_446_  (.A1(\soc/ram_ready ),
    .A2(\soc/_187_ ),
    .B1(\soc/_188_ ),
    .Y(\soc/_189_ ));
 sky130_fd_sc_hd__inv_1 \soc/_447_  (.A(\soc/spimem_rdata[23] ),
    .Y(\soc/_190_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_448_  (.A1(net110),
    .A2(\soc/_190_ ),
    .B1(\soc/_030_ ),
    .Y(\soc/_191_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_449_  (.A1(\iomem_rdata[23] ),
    .A2(\soc/_030_ ),
    .B1(\soc/_189_ ),
    .B2(\soc/_191_ ),
    .X(\soc/mem_rdata[23] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_450_  (.A1(\soc/simpleuart_reg_div_do[24] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net465),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_192_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_451_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[24] ),
    .B1(net112),
    .Y(\soc/_193_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_452_  (.A1(\soc/ram_ready ),
    .A2(\soc/_192_ ),
    .B1(\soc/_193_ ),
    .Y(\soc/_194_ ));
 sky130_fd_sc_hd__inv_1 \soc/_453_  (.A(\soc/spimem_rdata[24] ),
    .Y(\soc/_195_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_454_  (.A1(net110),
    .A2(\soc/_195_ ),
    .B1(net150),
    .Y(\soc/_196_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_455_  (.A1(\iomem_rdata[24] ),
    .A2(net150),
    .B1(\soc/_194_ ),
    .B2(\soc/_196_ ),
    .X(\soc/mem_rdata[24] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_456_  (.A1(\soc/simpleuart_reg_div_do[25] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net466),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_197_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_457_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[25] ),
    .B1(net112),
    .Y(\soc/_198_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_458_  (.A1(\soc/ram_ready ),
    .A2(\soc/_197_ ),
    .B1(\soc/_198_ ),
    .Y(\soc/_199_ ));
 sky130_fd_sc_hd__inv_1 \soc/_459_  (.A(\soc/spimem_rdata[25] ),
    .Y(\soc/_200_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_460_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_200_ ),
    .B1(net147),
    .Y(\soc/_201_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_461_  (.A1(net966),
    .A2(net148),
    .B1(\soc/_199_ ),
    .B2(\soc/_201_ ),
    .X(\soc/mem_rdata[25] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_462_  (.A1(\soc/simpleuart_reg_div_do[26] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net467),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_202_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_463_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[26] ),
    .B1(net112),
    .Y(\soc/_203_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_464_  (.A1(\soc/ram_ready ),
    .A2(\soc/_202_ ),
    .B1(\soc/_203_ ),
    .Y(\soc/_204_ ));
 sky130_fd_sc_hd__inv_1 \soc/_465_  (.A(\soc/spimem_rdata[26] ),
    .Y(\soc/_205_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_466_  (.A1(\soc/spimem_ready ),
    .A2(\soc/_205_ ),
    .B1(net148),
    .Y(\soc/_206_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_467_  (.A1(net868),
    .A2(net148),
    .B1(\soc/_204_ ),
    .B2(\soc/_206_ ),
    .X(\soc/mem_rdata[26] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_468_  (.A1(\soc/simpleuart_reg_div_do[27] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net468),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_207_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_469_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[27] ),
    .B1(net112),
    .Y(\soc/_208_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_470_  (.A1(\soc/ram_ready ),
    .A2(\soc/_207_ ),
    .B1(\soc/_208_ ),
    .Y(\soc/_209_ ));
 sky130_fd_sc_hd__inv_1 \soc/_471_  (.A(\soc/spimem_rdata[27] ),
    .Y(\soc/_210_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_472_  (.A1(net110),
    .A2(\soc/_210_ ),
    .B1(net148),
    .Y(\soc/_211_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_473_  (.A1(net787),
    .A2(net148),
    .B1(\soc/_209_ ),
    .B2(\soc/_211_ ),
    .X(\soc/mem_rdata[27] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_474_  (.A1(\soc/simpleuart_reg_div_do[28] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net469),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_212_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_475_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[28] ),
    .B1(net112),
    .Y(\soc/_213_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_476_  (.A1(\soc/ram_ready ),
    .A2(\soc/_212_ ),
    .B1(\soc/_213_ ),
    .Y(\soc/_214_ ));
 sky130_fd_sc_hd__inv_1 \soc/_477_  (.A(\soc/spimem_rdata[28] ),
    .Y(\soc/_215_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_478_  (.A1(net110),
    .A2(\soc/_215_ ),
    .B1(net150),
    .Y(\soc/_216_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_479_  (.A1(net833),
    .A2(net150),
    .B1(\soc/_214_ ),
    .B2(\soc/_216_ ),
    .X(\soc/mem_rdata[28] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_480_  (.A1(\soc/simpleuart_reg_div_do[29] ),
    .A2(\soc/_034_ ),
    .B1(net135),
    .B2(net470),
    .C1(\soc/_025_ ),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_217_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_481_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[29] ),
    .B1(net112),
    .Y(\soc/_218_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_482_  (.A1(\soc/ram_ready ),
    .A2(\soc/_217_ ),
    .B1(\soc/_218_ ),
    .Y(\soc/_219_ ));
 sky130_fd_sc_hd__inv_1 \soc/_483_  (.A(\soc/spimem_rdata[29] ),
    .Y(\soc/_220_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_484_  (.A1(net110),
    .A2(\soc/_220_ ),
    .B1(net150),
    .Y(\soc/_221_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_485_  (.A1(net816),
    .A2(net150),
    .B1(\soc/_219_ ),
    .B2(\soc/_221_ ),
    .X(\soc/mem_rdata[29] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_486_  (.A1(\soc/simpleuart_reg_div_do[30] ),
    .A2(net136),
    .B1(net134),
    .B2(net471),
    .C1(net138),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_222_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_487_  (.A1(net415),
    .A2(\soc/ram_rdata[30] ),
    .B1(net108),
    .Y(\soc/_223_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_488_  (.A1(net415),
    .A2(\soc/_222_ ),
    .B1(\soc/_223_ ),
    .Y(\soc/_224_ ));
 sky130_fd_sc_hd__inv_1 \soc/_489_  (.A(\soc/spimem_rdata[30] ),
    .Y(\soc/_225_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_490_  (.A1(net111),
    .A2(\soc/_225_ ),
    .B1(net146),
    .Y(\soc/_226_ ));
 sky130_fd_sc_hd__a22o_4 \soc/_491_  (.A1(\iomem_rdata[30] ),
    .A2(net146),
    .B1(\soc/_224_ ),
    .B2(\soc/_226_ ),
    .X(\soc/mem_rdata[30] ));
 sky130_fd_sc_hd__a222oi_1 \soc/_492_  (.A1(\soc/simpleuart_reg_div_do[31] ),
    .A2(net137),
    .B1(net135),
    .B2(\soc/spimemio/config_en ),
    .C1(net139),
    .C2(\soc/simpleuart_reg_dat_do[31] ),
    .Y(\soc/_227_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_493_  (.A1(\soc/ram_ready ),
    .A2(\soc/ram_rdata[31] ),
    .B1(net112),
    .Y(\soc/_228_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/_494_  (.A1(\soc/ram_ready ),
    .A2(\soc/_227_ ),
    .B1(\soc/_228_ ),
    .Y(\soc/_229_ ));
 sky130_fd_sc_hd__inv_1 \soc/_495_  (.A(\soc/spimem_rdata[31] ),
    .Y(\soc/_230_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/_496_  (.A1(net110),
    .A2(\soc/_230_ ),
    .B1(net148),
    .Y(\soc/_231_ ));
 sky130_fd_sc_hd__a22o_2 \soc/_497_  (.A1(net896),
    .A2(net148),
    .B1(\soc/_229_ ),
    .B2(\soc/_231_ ),
    .X(\soc/mem_rdata[31] ));
 sky130_fd_sc_hd__and2_0 \soc/_498_  (.A(net410),
    .B(net138),
    .X(\soc/_012_ ));
 sky130_fd_sc_hd__dfxtp_4 \soc/_499_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/_000_ ),
    .Q(\soc/ram_ready ));
 sky130_fd_sc_hd__conb_1 \soc/_243__448  (.LO(net448));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_04872_  (.A(\soc/cpu/latched_branch ),
    .B(\soc/cpu/irq_state[1] ),
    .C(\soc/cpu/irq_state[0] ),
    .Y(\soc/cpu/_00704_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04873_  (.A(\soc/cpu/prefetched_high_word ),
    .B(\soc/cpu/clear_prefetched_high_word_q ),
    .Y(\soc/cpu/_00705_ ));
 sky130_fd_sc_hd__nand3_2 \soc/cpu/_04874_  (.A(_074_),
    .B(\soc/cpu/_00704_ ),
    .C(\soc/cpu/_00705_ ),
    .Y(\soc/cpu/clear_prefetched_high_word ));
 sky130_fd_sc_hd__and2_4 \soc/cpu/_04876_  (.A(\soc/cpu/latched_store ),
    .B(\soc/cpu/latched_branch ),
    .X(\soc/cpu/_00707_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_04877_  (.A(\soc/cpu/reg_next_pc[1] ),
    .B(\soc/cpu/_00707_ ),
    .Y(\soc/cpu/_00708_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_04878_  (.A(\soc/cpu/latched_store ),
    .B(\soc/cpu/latched_branch ),
    .Y(\soc/cpu/_00709_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_04880_  (.A(\soc/cpu/mem_do_prefetch ),
    .B(\soc/cpu/mem_do_rinst ),
    .X(\soc/cpu/_00711_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_04881_  (.A1(\soc/cpu/reg_out[1] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_00711_ ),
    .Y(\soc/cpu/_00712_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_04882_  (.A(\soc/cpu/mem_la_secondword ),
    .B(\soc/cpu/_00708_ ),
    .C(\soc/cpu/_00712_ ),
    .Y(\soc/cpu/_00713_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04883_  (.A(\soc/cpu/prefetched_high_word ),
    .B(\soc/cpu/_00713_ ),
    .Y(\soc/cpu/_00714_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_04884_  (.A(\soc/cpu/clear_prefetched_high_word ),
    .B(\soc/cpu/_00714_ ),
    .Y(\soc/cpu/_00715_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_04885_  (.A(\soc/cpu/mem_la_secondword ),
    .B(\soc/cpu/_00715_ ),
    .Y(\soc/cpu/_00716_ ));
 sky130_fd_sc_hd__a22o_4 \soc/cpu/_04887_  (.A1(\soc/mem_valid ),
    .A2(\soc/mem_ready ),
    .B1(\soc/cpu/_00715_ ),
    .B2(\soc/cpu/mem_do_rinst ),
    .X(\soc/cpu/_00718_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_04890_  (.A1(\soc/mem_valid ),
    .A2(\soc/mem_ready ),
    .B1(\soc/cpu/_00715_ ),
    .B2(\soc/cpu/mem_do_rinst ),
    .Y(\soc/cpu/_00721_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04892_  (.A(\soc/cpu/mem_rdata_q[0] ),
    .B(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_00723_ ));
 sky130_fd_sc_hd__a21boi_1 \soc/cpu/_04893_  (.A1(\soc/mem_rdata[0] ),
    .A2(\soc/cpu/_00718_ ),
    .B1_N(\soc/cpu/_00723_ ),
    .Y(\soc/cpu/_00724_ ));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_04894_  (.A(\soc/cpu/mem_la_secondword ),
    .B(\soc/cpu/_00708_ ),
    .C(\soc/cpu/_00712_ ),
    .X(\soc/cpu/_00725_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_04896_  (.A0(\soc/mem_rdata[16] ),
    .A1(\soc/cpu/mem_rdata_q[16] ),
    .S(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_00727_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_04897_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_00727_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_00728_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_04898_  (.A1(\soc/cpu/_00713_ ),
    .A2(\soc/cpu/_00724_ ),
    .B1(\soc/cpu/_00728_ ),
    .Y(\soc/cpu/_00729_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_04899_  (.A1(\soc/cpu/mem_16bit_buffer[0] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_00729_ ),
    .X(\soc/cpu/_00730_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04901_  (.A(\soc/cpu/mem_rdata_q[1] ),
    .B(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_00732_ ));
 sky130_fd_sc_hd__a21boi_1 \soc/cpu/_04902_  (.A1(\soc/mem_rdata[1] ),
    .A2(\soc/cpu/_00718_ ),
    .B1_N(\soc/cpu/_00732_ ),
    .Y(\soc/cpu/_00733_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_04903_  (.A0(\soc/cpu/mem_rdata_q[17] ),
    .A1(\soc/mem_rdata[17] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_00734_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_04904_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_00734_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_00735_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_04905_  (.A1(\soc/cpu/_00713_ ),
    .A2(\soc/cpu/_00733_ ),
    .B1(\soc/cpu/_00735_ ),
    .Y(\soc/cpu/_00736_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_04906_  (.A1(\soc/cpu/mem_16bit_buffer[1] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_00736_ ),
    .X(\soc/cpu/_00737_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_04907_  (.A(\soc/cpu/_00730_ ),
    .B(\soc/cpu/_00737_ ),
    .Y(\soc/cpu/_00738_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04908_  (.A(\soc/cpu/mem_la_firstword_reg ),
    .B(\soc/cpu/last_mem_valid ),
    .Y(\soc/cpu/_00739_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_04909_  (.A1(\soc/cpu/last_mem_valid ),
    .A2(\soc/cpu/_00725_ ),
    .B1(\soc/cpu/_00739_ ),
    .Y(\soc/cpu/_00740_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_04910_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_00740_ ),
    .Y(\soc/cpu/_00741_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_04911_  (.A(\soc/cpu/mem_state[0] ),
    .B(\soc/cpu/mem_state[1] ),
    .Y(\soc/cpu/_00742_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_04912_  (.A1(\soc/cpu/mem_do_rdata ),
    .A2(\soc/cpu/_00711_ ),
    .B1(\soc/cpu/_00742_ ),
    .Y(\soc/cpu/_00743_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_04913_  (.A1(\soc/cpu/mem_la_secondword ),
    .A2(\soc/cpu/_00738_ ),
    .A3(\soc/cpu/_00741_ ),
    .B1(\soc/cpu/_00743_ ),
    .B2(\soc/cpu/_00715_ ),
    .Y(\soc/cpu/_00744_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04914_  (.A(_074_),
    .B(\soc/cpu/_00744_ ),
    .Y(\soc/cpu/_00745_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_04915_  (.A(\soc/cpu/_00745_ ),
    .Y(\soc/cpu/mem_la_read ));
 sky130_fd_sc_hd__inv_6 \soc/cpu/_04916_  (.A(\soc/cpu/decoder_trigger ),
    .Y(\soc/cpu/_00746_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04917_  (.A(\soc/cpu/irq_pending[29] ),
    .SLEEP(\soc/cpu/irq_mask[29] ),
    .X(\soc/cpu/_00747_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04918_  (.A(\soc/cpu/irq_pending[10] ),
    .SLEEP(\soc/cpu/irq_mask[10] ),
    .X(\soc/cpu/_00748_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04919_  (.A(\soc/cpu/irq_pending[20] ),
    .SLEEP(\soc/cpu/irq_mask[20] ),
    .X(\soc/cpu/_00749_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04920_  (.A(\soc/cpu/irq_pending[18] ),
    .SLEEP(net866),
    .X(\soc/cpu/_00750_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04921_  (.A(\soc/cpu/_00747_ ),
    .B(\soc/cpu/_00748_ ),
    .C(\soc/cpu/_00749_ ),
    .D(\soc/cpu/_00750_ ),
    .Y(\soc/cpu/_00751_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04922_  (.A(\soc/cpu/irq_pending[25] ),
    .SLEEP(\soc/cpu/irq_mask[25] ),
    .X(\soc/cpu/_00752_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04923_  (.A(\soc/cpu/irq_pending[1] ),
    .SLEEP(\soc/cpu/irq_mask[1] ),
    .X(\soc/cpu/_00753_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04924_  (.A(\soc/cpu/irq_pending[5] ),
    .SLEEP(\soc/cpu/irq_mask[5] ),
    .X(\soc/cpu/_00754_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04925_  (.A(\soc/cpu/irq_pending[12] ),
    .SLEEP(\soc/cpu/irq_mask[12] ),
    .X(\soc/cpu/_00755_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04926_  (.A(\soc/cpu/_00752_ ),
    .B(\soc/cpu/_00753_ ),
    .C(\soc/cpu/_00754_ ),
    .D(\soc/cpu/_00755_ ),
    .Y(\soc/cpu/_00756_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04927_  (.A(\soc/cpu/irq_pending[28] ),
    .SLEEP(\soc/cpu/irq_mask[28] ),
    .X(\soc/cpu/_00757_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_8 \soc/cpu/_04928_  (.A(\soc/cpu/irq_pending[7] ),
    .SLEEP(\soc/cpu/irq_mask[7] ),
    .X(\soc/cpu/_00758_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04929_  (.A(\soc/cpu/irq_pending[4] ),
    .SLEEP(\soc/cpu/irq_mask[4] ),
    .X(\soc/cpu/_00759_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04930_  (.A(\soc/cpu/irq_pending[27] ),
    .SLEEP(\soc/cpu/irq_mask[27] ),
    .X(\soc/cpu/_00760_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04931_  (.A(\soc/cpu/_00757_ ),
    .B(\soc/cpu/_00758_ ),
    .C(\soc/cpu/_00759_ ),
    .D(\soc/cpu/_00760_ ),
    .Y(\soc/cpu/_00761_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04932_  (.A(net856),
    .SLEEP(\soc/cpu/irq_mask[2] ),
    .X(\soc/cpu/_00762_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04933_  (.A(\soc/cpu/irq_pending[14] ),
    .SLEEP(\soc/cpu/irq_mask[14] ),
    .X(\soc/cpu/_00763_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04934_  (.A(\soc/cpu/irq_pending[21] ),
    .SLEEP(\soc/cpu/irq_mask[21] ),
    .X(\soc/cpu/_00764_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04935_  (.A(\soc/cpu/irq_pending[8] ),
    .SLEEP(\soc/cpu/irq_mask[8] ),
    .X(\soc/cpu/_00765_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04936_  (.A(\soc/cpu/_00762_ ),
    .B(\soc/cpu/_00763_ ),
    .C(\soc/cpu/_00764_ ),
    .D(\soc/cpu/_00765_ ),
    .Y(\soc/cpu/_00766_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_04937_  (.A(\soc/cpu/_00751_ ),
    .B(\soc/cpu/_00756_ ),
    .C(\soc/cpu/_00761_ ),
    .D(\soc/cpu/_00766_ ),
    .Y(\soc/cpu/_00767_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04938_  (.A(\soc/cpu/irq_pending[23] ),
    .SLEEP(\soc/cpu/irq_mask[23] ),
    .X(\soc/cpu/_00768_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04939_  (.A(\soc/cpu/irq_pending[30] ),
    .SLEEP(\soc/cpu/irq_mask[30] ),
    .X(\soc/cpu/_00769_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04940_  (.A(\soc/cpu/irq_pending[17] ),
    .SLEEP(\soc/cpu/irq_mask[17] ),
    .X(\soc/cpu/_00770_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04941_  (.A(\soc/cpu/irq_pending[3] ),
    .SLEEP(\soc/cpu/irq_mask[3] ),
    .X(\soc/cpu/_00771_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04942_  (.A(\soc/cpu/_00768_ ),
    .B(\soc/cpu/_00769_ ),
    .C(\soc/cpu/_00770_ ),
    .D(\soc/cpu/_00771_ ),
    .Y(\soc/cpu/_00772_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04943_  (.A(\soc/cpu/irq_pending[15] ),
    .SLEEP(\soc/cpu/irq_mask[15] ),
    .X(\soc/cpu/_00773_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04944_  (.A(\soc/cpu/irq_pending[9] ),
    .SLEEP(\soc/cpu/irq_mask[9] ),
    .X(\soc/cpu/_00774_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04945_  (.A(\soc/cpu/irq_pending[26] ),
    .SLEEP(\soc/cpu/irq_mask[26] ),
    .X(\soc/cpu/_00775_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04946_  (.A(\soc/cpu/irq_pending[6] ),
    .SLEEP(\soc/cpu/irq_mask[6] ),
    .X(\soc/cpu/_00776_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04947_  (.A(\soc/cpu/_00773_ ),
    .B(\soc/cpu/_00774_ ),
    .C(\soc/cpu/_00775_ ),
    .D(\soc/cpu/_00776_ ),
    .Y(\soc/cpu/_00777_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04948_  (.A(\soc/cpu/irq_pending[31] ),
    .SLEEP(\soc/cpu/irq_mask[31] ),
    .X(\soc/cpu/_00778_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04949_  (.A(\soc/cpu/irq_pending[19] ),
    .SLEEP(\soc/cpu/irq_mask[19] ),
    .X(\soc/cpu/_00779_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04950_  (.A(\soc/cpu/irq_pending[24] ),
    .SLEEP(\soc/cpu/irq_mask[24] ),
    .X(\soc/cpu/_00780_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04951_  (.A(\soc/cpu/irq_pending[16] ),
    .SLEEP(\soc/cpu/irq_mask[16] ),
    .X(\soc/cpu/_00781_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04952_  (.A(\soc/cpu/_00778_ ),
    .B(\soc/cpu/_00779_ ),
    .C(\soc/cpu/_00780_ ),
    .D(\soc/cpu/_00781_ ),
    .Y(\soc/cpu/_00782_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04953_  (.A(\soc/cpu/irq_pending[22] ),
    .SLEEP(\soc/cpu/irq_mask[22] ),
    .X(\soc/cpu/_00783_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04954_  (.A(\soc/cpu/irq_pending[11] ),
    .SLEEP(\soc/cpu/irq_mask[11] ),
    .X(\soc/cpu/_00784_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_04955_  (.A(\soc/cpu/irq_pending[0] ),
    .SLEEP(\soc/cpu/irq_mask[0] ),
    .X(\soc/cpu/_00785_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_04956_  (.A(\soc/cpu/irq_pending[13] ),
    .SLEEP(\soc/cpu/irq_mask[13] ),
    .X(\soc/cpu/_00786_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_04957_  (.A(\soc/cpu/_00783_ ),
    .B(\soc/cpu/_00784_ ),
    .C(\soc/cpu/_00785_ ),
    .D(\soc/cpu/_00786_ ),
    .Y(\soc/cpu/_00787_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_04958_  (.A(\soc/cpu/_00772_ ),
    .B(\soc/cpu/_00777_ ),
    .C(\soc/cpu/_00782_ ),
    .D(\soc/cpu/_00787_ ),
    .Y(\soc/cpu/_00788_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_04959_  (.A(\soc/cpu/_00767_ ),
    .B(\soc/cpu/_00788_ ),
    .Y(\soc/cpu/_00789_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_04960_  (.A(\soc/cpu/_00746_ ),
    .B(\soc/cpu/irq_active ),
    .C(\soc/cpu/irq_delay ),
    .D(\soc/cpu/_00789_ ),
    .Y(\soc/cpu/_00790_ ));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_04961_  (.A(\soc/cpu/irq_state[1] ),
    .B(\soc/cpu/irq_state[0] ),
    .C(\soc/cpu/_00790_ ),
    .X(\soc/cpu/_00791_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_04965_  (.A(_074_),
    .B(net819),
    .Y(\soc/cpu/_00795_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_04966_  (.A(\soc/cpu/_00791_ ),
    .B(\soc/cpu/_00795_ ),
    .Y(\soc/cpu/_00796_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_04967_  (.A1(\soc/cpu/decoder_trigger ),
    .A2(\soc/cpu/do_waitirq ),
    .B1(\soc/cpu/instr_waitirq ),
    .Y(\soc/cpu/_00797_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_04970_  (.A(\soc/cpu/mem_do_rinst ),
    .B(_074_),
    .C(\soc/cpu/reg_next_pc[0] ),
    .X(\soc/cpu/_00800_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_04971_  (.A(\soc/cpu/irq_active ),
    .B(\soc/cpu/irq_mask[2] ),
    .Y(\soc/cpu/_00801_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_04972_  (.A(\soc/cpu/_00800_ ),
    .B(\soc/cpu/_00801_ ),
    .Y(\soc/cpu/_00802_ ));
 sky130_fd_sc_hd__nand3_2 \soc/cpu/_04973_  (.A(\soc/cpu/mem_do_rinst ),
    .B(_074_),
    .C(\soc/cpu/reg_next_pc[0] ),
    .Y(\soc/cpu/_00803_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_04975_  (.A1(\soc/cpu/mem_do_rdata ),
    .A2(\soc/cpu/mem_do_wdata ),
    .B1(_074_),
    .Y(\soc/cpu/_00805_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_04976_  (.A(\soc/cpu/_00803_ ),
    .B(\soc/cpu/_00805_ ),
    .Y(\soc/cpu/_00806_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_04977_  (.A(\soc/cpu/irq_active ),
    .B(\soc/cpu/irq_mask[2] ),
    .C(\soc/cpu/_00800_ ),
    .D(\soc/cpu/_00805_ ),
    .Y(\soc/cpu/_00807_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04978_  (.A(\soc/cpu/pcpi_rs1 [0]),
    .B(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_00808_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_04981_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/pcpi_rs1 [1]),
    .B1(\soc/cpu/mem_wordsize[0] ),
    .Y(\soc/cpu/_00811_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_04982_  (.A(\soc/cpu/_00808_ ),
    .B(\soc/cpu/_00811_ ),
    .X(\soc/cpu/_00812_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04983_  (.A(\soc/cpu/_00803_ ),
    .B(\soc/cpu/_00812_ ),
    .Y(\soc/cpu/_00813_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_04984_  (.A(\soc/cpu/_00805_ ),
    .B(\soc/cpu/_00813_ ),
    .Y(\soc/cpu/_00814_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_04985_  (.A(\soc/cpu/_00807_ ),
    .B(\soc/cpu/_00814_ ),
    .Y(\soc/cpu/_00815_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_04986_  (.A(\soc/cpu/_00802_ ),
    .B(\soc/cpu/_00806_ ),
    .C(\soc/cpu/_00815_ ),
    .Y(\soc/cpu/_00816_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_04988_  (.A(\soc/cpu/instr_jal ),
    .B(\soc/cpu/_00746_ ),
    .Y(\soc/cpu/_00818_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_04989_  (.A(\soc/cpu/_00796_ ),
    .B(\soc/cpu/_00797_ ),
    .C(\soc/cpu/_00816_ ),
    .D(\soc/cpu/_00818_ ),
    .X(\soc/cpu/_00066_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_04993_  (.A(_074_),
    .B(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_00822_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_04996_  (.A1(\soc/cpu/mem_16bit_buffer[0] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_00729_ ),
    .Y(\soc/cpu/_00825_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_04997_  (.A1(\soc/cpu/mem_16bit_buffer[1] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_00736_ ),
    .Y(\soc/cpu/_00826_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_04998_  (.A(\soc/cpu/_00825_ ),
    .B(\soc/cpu/_00826_ ),
    .Y(\soc/cpu/_00827_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05000_  (.A1(net65),
    .A2(\soc/cpu/_00827_ ),
    .B1(\soc/cpu/_00713_ ),
    .Y(\soc/cpu/_00829_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05001_  (.A(\soc/cpu/mem_do_rinst ),
    .B(\soc/cpu/mem_do_rdata ),
    .C(\soc/cpu/mem_do_wdata ),
    .Y(\soc/cpu/_00830_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05002_  (.A(\soc/cpu/mem_do_rinst ),
    .B(\soc/cpu/mem_state[0] ),
    .C(\soc/cpu/mem_state[1] ),
    .Y(\soc/cpu/_00831_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_05003_  (.A1(\soc/cpu/_00742_ ),
    .A2(\soc/cpu/_00721_ ),
    .A3(\soc/cpu/_00830_ ),
    .B1(\soc/cpu/_00831_ ),
    .Y(\soc/cpu/_00832_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_05004_  (.A(_074_),
    .B(\soc/cpu/_00829_ ),
    .C(\soc/cpu/_00832_ ),
    .Y(\soc/cpu/_00833_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05005_  (.A1(net799),
    .A2(\soc/cpu/_00833_ ),
    .B1(\soc/cpu/mem_do_rdata ),
    .Y(\soc/cpu/_00834_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_05006_  (.A(\soc/cpu/instr_lh ),
    .B(\soc/cpu/instr_lhu ),
    .C(\soc/cpu/instr_lb ),
    .D(\soc/cpu/instr_lbu ),
    .X(\soc/cpu/_00835_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05007_  (.A(\soc/cpu/instr_lw ),
    .B(\soc/cpu/_00835_ ),
    .Y(\soc/cpu/_00836_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05008_  (.A(\soc/cpu/mem_do_rdata ),
    .B(\soc/cpu/_00822_ ),
    .Y(\soc/cpu/_00837_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_05009_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/cpu_state[5] ),
    .Y(\soc/cpu/_00838_ ));
 sky130_fd_sc_hd__inv_16 \soc/cpu/_05010_  (.A(\soc/cpu/cpu_state[1] ),
    .Y(\soc/cpu/_00839_ ));
 sky130_fd_sc_hd__clkinv_16 \soc/cpu/_05011_  (.A(_074_),
    .Y(\soc/cpu/_00840_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_05012_  (.A1(\soc/cpu/_00836_ ),
    .A2(\soc/cpu/_00837_ ),
    .B1(\soc/cpu/_00838_ ),
    .B2(\soc/cpu/_00839_ ),
    .C1(net132),
    .Y(\soc/cpu/_00841_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05013_  (.A(\soc/cpu/mem_do_prefetch ),
    .B(\soc/cpu/_00833_ ),
    .Y(\soc/cpu/_00842_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05014_  (.A_N(\soc/cpu/mem_do_wdata ),
    .B(\soc/cpu/_00842_ ),
    .Y(\soc/cpu/_00843_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05015_  (.A(\soc/cpu/instr_sh ),
    .B(\soc/cpu/instr_sb ),
    .C(\soc/cpu/instr_sw ),
    .Y(\soc/cpu/_00844_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05016_  (.A(_074_),
    .B(\soc/cpu/cpu_state[5] ),
    .Y(\soc/cpu/_00845_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_05017_  (.A1(\soc/cpu/_00843_ ),
    .A2(\soc/cpu/_00844_ ),
    .B1_N(\soc/cpu/_00845_ ),
    .Y(\soc/cpu/_00846_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_05018_  (.A1(\soc/cpu/_00822_ ),
    .A2(\soc/cpu/_00834_ ),
    .B1(\soc/cpu/_00841_ ),
    .C1(\soc/cpu/_00846_ ),
    .Y(\soc/cpu/_00847_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05019_  (.A(\soc/cpu/mem_wordsize[2] ),
    .B(\soc/cpu/_00847_ ),
    .Y(\soc/cpu/_00848_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05020_  (.A(\soc/cpu/_00845_ ),
    .B(\soc/cpu/_00843_ ),
    .Y(\soc/cpu/_00849_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05021_  (.A(\soc/cpu/instr_sh ),
    .B(\soc/cpu/_00849_ ),
    .Y(\soc/cpu/_00850_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05022_  (.A(net800),
    .B(\soc/cpu/_00837_ ),
    .X(\soc/cpu/_00851_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05023_  (.A1(\soc/cpu/instr_lh ),
    .A2(\soc/cpu/instr_lhu ),
    .B1(\soc/cpu/_00851_ ),
    .Y(\soc/cpu/_00852_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05024_  (.A(\soc/cpu/_00848_ ),
    .B(\soc/cpu/_00850_ ),
    .C(\soc/cpu/_00852_ ),
    .Y(\soc/cpu/_00073_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05025_  (.A1(\soc/cpu/instr_lb ),
    .A2(\soc/cpu/instr_lbu ),
    .B1(\soc/cpu/_00851_ ),
    .Y(\soc/cpu/_00853_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_05028_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_00847_ ),
    .B1(\soc/cpu/_00849_ ),
    .B2(\soc/cpu/instr_sb ),
    .Y(\soc/cpu/_00856_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05029_  (.A(\soc/cpu/_00853_ ),
    .B(\soc/cpu/_00856_ ),
    .Y(\soc/cpu/_00072_ ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_05030_  (.A(_074_),
    .B(\soc/cpu/mem_do_wdata ),
    .C(\soc/cpu/_00742_ ),
    .X(\soc/cpu/_00857_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05032_  (.A(\soc/cpu/mem_wordsize[0] ),
    .B(\soc/cpu/_00847_ ),
    .Y(\soc/cpu/_00858_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_05033_  (.A(net132),
    .B(\soc/cpu/_00839_ ),
    .Y(\soc/cpu/_00859_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_05035_  (.A1(\soc/cpu/instr_sw ),
    .A2(\soc/cpu/_00849_ ),
    .B1(\soc/cpu/_00851_ ),
    .B2(\soc/cpu/instr_lw ),
    .C1(\soc/cpu/_00859_ ),
    .Y(\soc/cpu/_00861_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05036_  (.A(\soc/cpu/_00858_ ),
    .B(\soc/cpu/_00861_ ),
    .Y(\soc/cpu/_00071_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05038_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/mem_wordsize[2] ),
    .B1(\soc/cpu/_00811_ ),
    .Y(\soc/cpu/_00863_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05039_  (.A(\soc/cpu/_00807_ ),
    .B(\soc/cpu/_00863_ ),
    .Y(\soc/cpu/_00864_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05040_  (.A(\soc/cpu/_00802_ ),
    .B(\soc/cpu/_00864_ ),
    .Y(\soc/cpu/_00865_ ));
 sky130_fd_sc_hd__a32oi_2 \soc/cpu/_05041_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/mem_wordsize[2] ),
    .A3(\soc/cpu/_00807_ ),
    .B1(\soc/cpu/_00805_ ),
    .B2(\soc/cpu/_00803_ ),
    .Y(\soc/cpu/_00866_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05042_  (.A(\soc/cpu/_00813_ ),
    .B(\soc/cpu/_00866_ ),
    .Y(\soc/cpu/_00867_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05043_  (.A(\soc/cpu/_00865_ ),
    .B(\soc/cpu/_00867_ ),
    .Y(\soc/cpu/_00868_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_05047_  (.A(\soc/cpu/instr_maskirq ),
    .B(\soc/cpu/instr_retirq ),
    .C(\soc/cpu/instr_timer ),
    .Y(\soc/cpu/_00872_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_05048_  (.A(\soc/cpu/instr_rdinstrh ),
    .B(\soc/cpu/instr_rdinstr ),
    .C(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_00873_ ));
 sky130_fd_sc_hd__and2_4 \soc/cpu/_05049_  (.A(net160),
    .B(\soc/cpu/_00873_ ),
    .X(\soc/cpu/_00874_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_05050_  (.A(\soc/cpu/instr_waitirq ),
    .B(\soc/cpu/instr_fence ),
    .C(\soc/cpu/instr_and ),
    .D(\soc/cpu/instr_rdcycle ),
    .X(\soc/cpu/_00875_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05051_  (.A(\soc/cpu/instr_bgeu ),
    .B(\soc/cpu/instr_bge ),
    .C(\soc/cpu/_00875_ ),
    .Y(\soc/cpu/_00876_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05052_  (.A(\soc/cpu/instr_beq ),
    .B(\soc/cpu/instr_bne ),
    .C(\soc/cpu/instr_jalr ),
    .Y(\soc/cpu/_00877_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_05053_  (.A(\soc/cpu/instr_auipc ),
    .B(\soc/cpu/instr_lui ),
    .X(\soc/cpu/_00878_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05054_  (.A(\soc/cpu/instr_jal ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_00879_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05055_  (.A(net802),
    .B(\soc/cpu/instr_slt ),
    .C(net751),
    .D(\soc/cpu/instr_slti ),
    .Y(\soc/cpu/_00880_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05056_  (.A(\soc/cpu/_00844_ ),
    .B(\soc/cpu/_00877_ ),
    .C(\soc/cpu/_00879_ ),
    .D(\soc/cpu/_00880_ ),
    .Y(\soc/cpu/_00881_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05060_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/instr_sll ),
    .C(\soc/cpu/instr_srai ),
    .D(\soc/cpu/instr_add ),
    .Y(\soc/cpu/_00885_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05061_  (.A(\soc/cpu/instr_sra ),
    .B(\soc/cpu/instr_or ),
    .C(\soc/cpu/instr_xor ),
    .D(\soc/cpu/instr_srl ),
    .Y(\soc/cpu/_00886_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05062_  (.A(\soc/cpu/instr_xori ),
    .B(\soc/cpu/instr_addi ),
    .C(\soc/cpu/instr_bltu ),
    .D(\soc/cpu/instr_blt ),
    .Y(\soc/cpu/_00887_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05063_  (.A(\soc/cpu/instr_slli ),
    .B(\soc/cpu/instr_srli ),
    .C(\soc/cpu/instr_ori ),
    .D(\soc/cpu/instr_andi ),
    .Y(\soc/cpu/_00888_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05064_  (.A(\soc/cpu/_00885_ ),
    .B(\soc/cpu/_00886_ ),
    .C(\soc/cpu/_00887_ ),
    .D(\soc/cpu/_00888_ ),
    .Y(\soc/cpu/_00889_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05065_  (.A(\soc/cpu/_00881_ ),
    .B(\soc/cpu/_00889_ ),
    .Y(\soc/cpu/_00890_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_05066_  (.A(\soc/cpu/_00836_ ),
    .B(\soc/cpu/_00874_ ),
    .C(\soc/cpu/_00876_ ),
    .D(\soc/cpu/_00890_ ),
    .Y(\soc/cpu/_00891_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05067_  (.A(net953),
    .B(\soc/cpu/_00891_ ),
    .Y(\soc/cpu/_00892_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05069_  (.A(_074_),
    .B(\soc/cpu/cpu_state[2] ),
    .Y(\soc/cpu/_00894_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05074_  (.A(net799),
    .B(\soc/cpu/_00833_ ),
    .Y(\soc/cpu/_00899_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05075_  (.A(\soc/cpu/_00868_ ),
    .B(\soc/cpu/_00899_ ),
    .Y(\soc/cpu/_00900_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05076_  (.A(_074_),
    .B(\soc/cpu/cpu_state[6] ),
    .C(\soc/cpu/_00900_ ),
    .Y(\soc/cpu/_00901_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_05077_  (.A1(\soc/cpu/_00868_ ),
    .A2(\soc/cpu/_00892_ ),
    .A3(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_00901_ ),
    .Y(\soc/cpu/_00070_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05078_  (.A(\soc/cpu/mem_do_rdata ),
    .B(\soc/cpu/mem_do_wdata ),
    .Y(\soc/cpu/_00902_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05079_  (.A(\soc/cpu/_00800_ ),
    .B(\soc/cpu/_00801_ ),
    .C(\soc/cpu/_00902_ ),
    .D(\soc/cpu/_00812_ ),
    .Y(\soc/cpu/_00903_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05080_  (.A(\soc/cpu/irq_active ),
    .B(\soc/cpu/irq_mask[1] ),
    .Y(\soc/cpu/_00904_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05081_  (.A(\soc/cpu/_00891_ ),
    .Y(\soc/cpu/_00905_ ));
 sky130_fd_sc_hd__and2_4 \soc/cpu/_05082_  (.A(_074_),
    .B(net801),
    .X(\soc/cpu/_00906_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05084_  (.A(\soc/cpu/_00905_ ),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_00908_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_05085_  (.A1(\soc/cpu/_00803_ ),
    .A2(\soc/cpu/_00801_ ),
    .B1(\soc/cpu/_00904_ ),
    .B2(\soc/cpu/_00908_ ),
    .X(\soc/cpu/_00909_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05086_  (.A(\soc/cpu/_00802_ ),
    .B(\soc/cpu/_00815_ ),
    .Y(\soc/cpu/_00910_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05087_  (.A(\soc/cpu/cpu_state[0] ),
    .B(\soc/cpu/_00910_ ),
    .Y(\soc/cpu/_00911_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_05088_  (.A(\soc/cpu/cpu_state[0] ),
    .B(\soc/cpu/_00803_ ),
    .C(\soc/cpu/_00902_ ),
    .X(\soc/cpu/_00912_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05090_  (.A1(\soc/cpu/_00903_ ),
    .A2(\soc/cpu/_00912_ ),
    .B1(_074_),
    .Y(\soc/cpu/_00914_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_05091_  (.A1(\soc/cpu/_00903_ ),
    .A2(\soc/cpu/_00909_ ),
    .B1(\soc/cpu/_00911_ ),
    .C1(\soc/cpu/_00914_ ),
    .Y(\soc/cpu/_00064_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05094_  (.A(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .B(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_00917_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05095_  (.A1(\soc/cpu/mem_do_prefetch ),
    .A2(\soc/cpu/_00838_ ),
    .B1(\soc/cpu/_00917_ ),
    .Y(\soc/cpu/_00918_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05096_  (.A(\soc/cpu/_00816_ ),
    .B(\soc/cpu/_00918_ ),
    .Y(\soc/cpu/_00919_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05098_  (.A(\soc/cpu/_00806_ ),
    .B(\soc/cpu/_00815_ ),
    .Y(\soc/cpu/_00921_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05100_  (.A(\soc/cpu/decoder_trigger ),
    .B(\soc/cpu/do_waitirq ),
    .Y(\soc/cpu/_00923_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_05101_  (.A(\soc/cpu/instr_waitirq ),
    .SLEEP(\soc/cpu/_00923_ ),
    .X(\soc/cpu/_00924_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05102_  (.A(\soc/cpu/decoder_trigger ),
    .B(\soc/cpu/_00924_ ),
    .Y(\soc/cpu/_00925_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05103_  (.A(\soc/cpu/instr_jal ),
    .B(\soc/cpu/decoder_trigger ),
    .Y(\soc/cpu/_00926_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_05105_  (.A(\soc/cpu/_00746_ ),
    .B(\soc/cpu/instr_waitirq ),
    .Y(\soc/cpu/_00928_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_05106_  (.A1(\soc/cpu/_00924_ ),
    .A2(\soc/cpu/_00868_ ),
    .A3(\soc/cpu/_00926_ ),
    .B1(\soc/cpu/_00928_ ),
    .B2(\soc/cpu/_00802_ ),
    .Y(\soc/cpu/_00929_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05107_  (.A(\soc/cpu/_00797_ ),
    .B(\soc/cpu/_00815_ ),
    .Y(\soc/cpu/_00930_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05108_  (.A1(\soc/cpu/_00921_ ),
    .A2(\soc/cpu/_00925_ ),
    .B1(\soc/cpu/_00929_ ),
    .C1(\soc/cpu/_00930_ ),
    .Y(\soc/cpu/_00931_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05109_  (.A1(\soc/cpu/_00797_ ),
    .A2(\soc/cpu/_00806_ ),
    .B1(\soc/cpu/_00931_ ),
    .B2(\soc/cpu/_00791_ ),
    .Y(\soc/cpu/_00932_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05110_  (.A(\soc/cpu/cpu_state[1] ),
    .B(\soc/cpu/_00932_ ),
    .Y(\soc/cpu/_00933_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05111_  (.A(\soc/cpu/cpu_state[2] ),
    .B(\soc/cpu/_00905_ ),
    .Y(\soc/cpu/_00934_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05112_  (.A(\soc/cpu/irq_active ),
    .B(\soc/cpu/irq_mask[1] ),
    .C(\soc/cpu/_00934_ ),
    .Y(\soc/cpu/_00935_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_05113_  (.A(\soc/cpu/reg_sh[4] ),
    .B(\soc/cpu/reg_sh[2] ),
    .C(\soc/cpu/reg_sh[3] ),
    .Y(\soc/cpu/_00936_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05114_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/_00936_ ),
    .Y(\soc/cpu/_00937_ ));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_05115_  (.A(net804),
    .B(\soc/cpu/reg_sh[1] ),
    .C(\soc/cpu/_00937_ ),
    .X(\soc/cpu/_00938_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05116_  (.A_N(\soc/cpu/_00938_ ),
    .B(\soc/cpu/_00921_ ),
    .Y(\soc/cpu/_00939_ ));
 sky130_fd_sc_hd__clkinv_4 \soc/cpu/_05117_  (.A(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_00940_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05118_  (.A(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .B(\soc/cpu/_00940_ ),
    .Y(\soc/cpu/_00941_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05119_  (.A(\soc/cpu/_00867_ ),
    .B(\soc/cpu/_00941_ ),
    .Y(\soc/cpu/_00942_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05120_  (.A(\soc/cpu/_00865_ ),
    .B(\soc/cpu/_00941_ ),
    .Y(\soc/cpu/_00943_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05121_  (.A(_074_),
    .B(\soc/cpu/_00939_ ),
    .C(\soc/cpu/_00942_ ),
    .D(\soc/cpu/_00943_ ),
    .Y(\soc/cpu/_00944_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05122_  (.A(net160),
    .B(\soc/cpu/_00873_ ),
    .Y(\soc/cpu/_00945_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05123_  (.A(\soc/cpu/instr_rdcycle ),
    .B(\soc/cpu/_00945_ ),
    .Y(\soc/cpu/_00946_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05124_  (.A1(\soc/cpu/_00807_ ),
    .A2(\soc/cpu/_00863_ ),
    .B1(\soc/cpu/_00814_ ),
    .Y(\soc/cpu/_00947_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05125_  (.A(\soc/cpu/_00802_ ),
    .B(\soc/cpu/_00866_ ),
    .Y(\soc/cpu/_00948_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \soc/cpu/_05127_  (.A1_N(\soc/cpu/_00947_ ),
    .A2_N(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_00948_ ),
    .B2(\soc/cpu/cpu_state[2] ),
    .Y(\soc/cpu/_00950_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05128_  (.A(\soc/cpu/_00946_ ),
    .B(\soc/cpu/_00950_ ),
    .Y(\soc/cpu/_00951_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05129_  (.A1(\soc/cpu/irq_mask[1] ),
    .A2(\soc/cpu/_00908_ ),
    .B1(\soc/cpu/_00938_ ),
    .X(\soc/cpu/_00952_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05130_  (.A(net819),
    .B(\soc/cpu/_00791_ ),
    .Y(\soc/cpu/_00953_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05131_  (.A1(\soc/cpu/_00802_ ),
    .A2(\soc/cpu/_00952_ ),
    .B1(\soc/cpu/_00953_ ),
    .B2(\soc/cpu/_00868_ ),
    .Y(\soc/cpu/_00954_ ));
 sky130_fd_sc_hd__a2111oi_0 \soc/cpu/_05132_  (.A1(\soc/cpu/_00921_ ),
    .A2(\soc/cpu/_00935_ ),
    .B1(\soc/cpu/_00944_ ),
    .C1(\soc/cpu/_00951_ ),
    .D1(\soc/cpu/_00954_ ),
    .Y(\soc/cpu/_00955_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_05133_  (.A1(\soc/cpu/_00833_ ),
    .A2(\soc/cpu/_00919_ ),
    .B1(\soc/cpu/_00933_ ),
    .C1(\soc/cpu/_00955_ ),
    .Y(\soc/cpu/_00065_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05134_  (.A(_074_),
    .B(\soc/cpu/cpu_state[5] ),
    .C(\soc/cpu/_00900_ ),
    .Y(\soc/cpu/_00956_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05135_  (.A(\soc/cpu/is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .B(\soc/cpu/is_lui_auipc_jal ),
    .Y(\soc/cpu/_00957_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_05136_  (.A(\soc/cpu/_00892_ ),
    .B(\soc/cpu/_00946_ ),
    .C(\soc/cpu/_00957_ ),
    .X(\soc/cpu/_00958_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05138_  (.A(\soc/cpu/is_slli_srli_srai ),
    .B(\soc/cpu/_00868_ ),
    .C(\soc/cpu/_00905_ ),
    .D(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_00960_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05139_  (.A(net952),
    .B(\soc/cpu/_00958_ ),
    .C(\soc/cpu/_00960_ ),
    .Y(\soc/cpu/_00961_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05140_  (.A(\soc/cpu/_00956_ ),
    .B(\soc/cpu/_00961_ ),
    .Y(\soc/cpu/_00069_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05141_  (.A(\soc/cpu/_00879_ ),
    .Y(\soc/cpu/_00033_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_05142_  (.A(\soc/cpu/instr_slt ),
    .B(\soc/cpu/instr_slti ),
    .C(\soc/cpu/instr_blt ),
    .X(\soc/cpu/_00034_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_05143_  (.A(\soc/cpu/instr_sltu ),
    .B(net751),
    .C(\soc/cpu/instr_bltu ),
    .X(\soc/cpu/_00035_ ));
 sky130_fd_sc_hd__inv_4 \soc/cpu/_05145_  (.A(\soc/cpu/_00833_ ),
    .Y(\soc/cpu/_00963_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05146_  (.A(net132),
    .B(\soc/cpu/_00963_ ),
    .Y(\soc/cpu/_00964_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05147_  (.A(net954),
    .B(\soc/cpu/cpu_state[3] ),
    .C(\soc/cpu/_00816_ ),
    .D(\soc/cpu/_00964_ ),
    .Y(\soc/cpu/_00965_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_05148_  (.A(\soc/cpu/is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .B(\soc/cpu/is_lui_auipc_jal ),
    .X(\soc/cpu/_00966_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05151_  (.A(\soc/cpu/_00816_ ),
    .B(\soc/cpu/_00906_ ),
    .C(\soc/cpu/_00966_ ),
    .Y(\soc/cpu/_00969_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05153_  (.A(\soc/cpu/is_slli_srli_srai ),
    .B(net952),
    .C(\soc/cpu/_00868_ ),
    .Y(\soc/cpu/_00971_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05154_  (.A(_074_),
    .B(\soc/cpu/_00891_ ),
    .Y(\soc/cpu/_00972_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05155_  (.A(\soc/cpu/is_sll_srl_sra ),
    .B(\soc/cpu/_00972_ ),
    .Y(\soc/cpu/_00973_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05156_  (.A(net801),
    .B(\soc/cpu/_00958_ ),
    .C(\soc/cpu/_00971_ ),
    .D(\soc/cpu/_00973_ ),
    .Y(\soc/cpu/_00974_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05157_  (.A(\soc/cpu/_00965_ ),
    .B(\soc/cpu/_00969_ ),
    .C(\soc/cpu/_00974_ ),
    .Y(\soc/cpu/_00067_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05159_  (.A_N(net804),
    .B(\soc/cpu/_00936_ ),
    .Y(\soc/cpu/_00976_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/_05162_  (.A1(\soc/cpu/reg_sh[1] ),
    .A2(\soc/cpu/_00976_ ),
    .B1(\soc/cpu/cpu_state[4] ),
    .X(\soc/cpu/_00979_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05163_  (.A(\soc/cpu/_00816_ ),
    .B(\soc/cpu/_00958_ ),
    .Y(\soc/cpu/_00980_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05164_  (.A(net801),
    .B(\soc/cpu/is_sll_srl_sra ),
    .C(\soc/cpu/_00891_ ),
    .Y(\soc/cpu/_00981_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05165_  (.A(\soc/cpu/is_slli_srli_srai ),
    .B(\soc/cpu/_00980_ ),
    .C(\soc/cpu/_00981_ ),
    .Y(\soc/cpu/_00982_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05166_  (.A1(\soc/cpu/_00816_ ),
    .A2(\soc/cpu/_00979_ ),
    .B1(\soc/cpu/_00982_ ),
    .Y(\soc/cpu/_00983_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05167_  (.A(\soc/cpu/is_slli_srli_srai ),
    .B(\soc/cpu/_00816_ ),
    .C(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_00984_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05168_  (.A1(net131),
    .A2(\soc/cpu/_00983_ ),
    .B1(\soc/cpu/_00984_ ),
    .Y(\soc/cpu/_00068_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05169_  (.A(\soc/cpu/latched_store ),
    .Y(\soc/cpu/_00985_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_05170_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/cpuregs_waddr[0] ),
    .C(\soc/cpu/cpuregs_waddr[2] ),
    .D(\soc/cpu/cpuregs_waddr[4] ),
    .X(\soc/cpu/_00986_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05171_  (.A1(\soc/cpu/cpuregs_waddr[3] ),
    .A2(\soc/cpu/_00986_ ),
    .B1(\soc/cpu/_00859_ ),
    .Y(\soc/cpu/_00987_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_05172_  (.A1(\soc/cpu/_00985_ ),
    .A2(\soc/cpu/_00704_ ),
    .B1(\soc/cpu/_00987_ ),
    .Y(\soc/cpu/_00074_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_05174_  (.A(\soc/cpu/cpu_state[2] ),
    .B(\soc/cpu/cpu_state[4] ),
    .Y(\soc/cpu/_00989_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05175_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_00989_ ),
    .Y(\soc/cpu/_00990_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05176_  (.A(net778),
    .B(\soc/cpu/_00990_ ),
    .Y(\soc/cpu/_00991_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_05177_  (.A(\soc/cpu/irq_state[1] ),
    .B(\soc/cpu/_00940_ ),
    .C(\soc/cpu/_00991_ ),
    .Y(\soc/cpu/_00992_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_05180_  (.A1(\soc/cpu/irq_mask[2] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(_074_),
    .C1(\soc/cpu/irq_pending[2] ),
    .Y(\soc/cpu/_00995_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05181_  (.A(\soc/cpu/_00808_ ),
    .B(\soc/cpu/_00811_ ),
    .Y(\soc/cpu/_00996_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05182_  (.A1(\soc/cpu/_00807_ ),
    .A2(\soc/cpu/_00996_ ),
    .B1(net446),
    .Y(\soc/cpu/_00997_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05183_  (.A(\soc/cpu/_00802_ ),
    .B(\soc/cpu/_00995_ ),
    .C(\soc/cpu/_00997_ ),
    .Y(\soc/cpu/_00023_ ));
 sky130_fd_sc_hd__or3_2 \soc/cpu/_05184_  (.A(\soc/cpu/timer[1] ),
    .B(\soc/cpu/timer[0] ),
    .C(\soc/cpu/timer[2] ),
    .X(\soc/cpu/_00998_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05185_  (.A(\soc/cpu/timer[5] ),
    .B(\soc/cpu/timer[4] ),
    .C(\soc/cpu/timer[3] ),
    .D(\soc/cpu/_00998_ ),
    .Y(\soc/cpu/_00999_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_05186_  (.A(\soc/cpu/_00999_ ),
    .SLEEP(\soc/cpu/timer[6] ),
    .X(\soc/cpu/_01000_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_05187_  (.A_N(\soc/cpu/timer[7] ),
    .B(\soc/cpu/_01000_ ),
    .Y(\soc/cpu/_01001_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05188_  (.A(\soc/cpu/timer[9] ),
    .B(\soc/cpu/timer[8] ),
    .C(\soc/cpu/_01001_ ),
    .Y(\soc/cpu/_01002_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05189_  (.A_N(\soc/cpu/timer[10] ),
    .B(\soc/cpu/_01002_ ),
    .Y(\soc/cpu/_01003_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05190_  (.A(\soc/cpu/timer[11] ),
    .B(\soc/cpu/timer[12] ),
    .C(\soc/cpu/_01003_ ),
    .Y(\soc/cpu/_01004_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05191_  (.A_N(\soc/cpu/timer[13] ),
    .B(\soc/cpu/_01004_ ),
    .Y(\soc/cpu/_01005_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05192_  (.A(\soc/cpu/timer[15] ),
    .B(\soc/cpu/timer[14] ),
    .C(\soc/cpu/_01005_ ),
    .Y(\soc/cpu/_01006_ ));
 sky130_fd_sc_hd__nand2b_2 \soc/cpu/_05193_  (.A_N(\soc/cpu/timer[16] ),
    .B(\soc/cpu/_01006_ ),
    .Y(\soc/cpu/_01007_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05194_  (.A(\soc/cpu/timer[17] ),
    .B(\soc/cpu/timer[19] ),
    .C(\soc/cpu/timer[18] ),
    .D(\soc/cpu/_01007_ ),
    .Y(\soc/cpu/_01008_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05195_  (.A(\soc/cpu/timer[21] ),
    .B(\soc/cpu/timer[20] ),
    .Y(\soc/cpu/_01009_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05196_  (.A(\soc/cpu/_01008_ ),
    .B(\soc/cpu/_01009_ ),
    .Y(\soc/cpu/_01010_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05197_  (.A(\soc/cpu/timer[23] ),
    .B(\soc/cpu/timer[22] ),
    .C(\soc/cpu/_01010_ ),
    .Y(\soc/cpu/_01011_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05198_  (.A_N(\soc/cpu/timer[24] ),
    .B(\soc/cpu/_01011_ ),
    .Y(\soc/cpu/_01012_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05199_  (.A(\soc/cpu/timer[25] ),
    .B(\soc/cpu/timer[26] ),
    .C(\soc/cpu/_01012_ ),
    .Y(\soc/cpu/_01013_ ));
 sky130_fd_sc_hd__nand2b_2 \soc/cpu/_05200_  (.A_N(\soc/cpu/timer[27] ),
    .B(\soc/cpu/_01013_ ),
    .Y(\soc/cpu/_01014_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05201_  (.A(\soc/cpu/timer[28] ),
    .B(\soc/cpu/_01014_ ),
    .Y(\soc/cpu/_01015_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05202_  (.A(\soc/cpu/timer[29] ),
    .B(\soc/cpu/_01015_ ),
    .Y(\soc/cpu/_01016_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05203_  (.A1(\soc/cpu/timer[25] ),
    .A2(\soc/cpu/_01012_ ),
    .B1(\soc/cpu/timer[26] ),
    .X(\soc/cpu/_01017_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05204_  (.A(\soc/cpu/_01013_ ),
    .B(\soc/cpu/_01017_ ),
    .Y(\soc/cpu/_01018_ ));
 sky130_fd_sc_hd__xor2_2 \soc/cpu/_05205_  (.A(\soc/cpu/timer[22] ),
    .B(\soc/cpu/_01010_ ),
    .X(\soc/cpu/_01019_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05206_  (.A(\soc/cpu/timer[17] ),
    .B(\soc/cpu/timer[18] ),
    .C(\soc/cpu/_01007_ ),
    .Y(\soc/cpu/_01020_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05207_  (.A(\soc/cpu/timer[19] ),
    .B(\soc/cpu/_01020_ ),
    .Y(\soc/cpu/_01021_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05208_  (.A(\soc/cpu/timer[14] ),
    .B(\soc/cpu/_01005_ ),
    .Y(\soc/cpu/_01022_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05209_  (.A(\soc/cpu/timer[11] ),
    .B(\soc/cpu/_01003_ ),
    .X(\soc/cpu/_01023_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05210_  (.A1(\soc/cpu/timer[8] ),
    .A2(\soc/cpu/_01001_ ),
    .B1(\soc/cpu/timer[9] ),
    .X(\soc/cpu/_01024_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05211_  (.A(\soc/cpu/_01002_ ),
    .B(\soc/cpu/_01024_ ),
    .Y(\soc/cpu/_01025_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05212_  (.A(\soc/cpu/timer[8] ),
    .B(\soc/cpu/_01001_ ),
    .X(\soc/cpu/_01026_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05213_  (.A(\soc/cpu/timer[6] ),
    .B(\soc/cpu/_00999_ ),
    .Y(\soc/cpu/_01027_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05214_  (.A(\soc/cpu/timer[4] ),
    .B(\soc/cpu/timer[3] ),
    .C(\soc/cpu/_00998_ ),
    .Y(\soc/cpu/_01028_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05215_  (.A(\soc/cpu/timer[5] ),
    .B(\soc/cpu/_01028_ ),
    .Y(\soc/cpu/_01029_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05216_  (.A(\soc/cpu/timer[3] ),
    .B(\soc/cpu/timer[2] ),
    .C(\soc/cpu/timer[17] ),
    .D(\soc/cpu/timer[18] ),
    .Y(\soc/cpu/_01030_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05217_  (.A(\soc/cpu/_01009_ ),
    .B(\soc/cpu/_01030_ ),
    .Y(\soc/cpu/_01031_ ));
 sky130_fd_sc_hd__nor4b_1 \soc/cpu/_05218_  (.A(\soc/cpu/timer[4] ),
    .B(\soc/cpu/timer[7] ),
    .C(\soc/cpu/timer[1] ),
    .D_N(\soc/cpu/timer[0] ),
    .Y(\soc/cpu/_01032_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05219_  (.A(\soc/cpu/timer[10] ),
    .B(\soc/cpu/timer[13] ),
    .C(\soc/cpu/timer[12] ),
    .D(\soc/cpu/timer[15] ),
    .Y(\soc/cpu/_01033_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05220_  (.A(\soc/cpu/timer[28] ),
    .B(\soc/cpu/timer[31] ),
    .C(\soc/cpu/timer[30] ),
    .Y(\soc/cpu/_01034_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05221_  (.A(\soc/cpu/timer[23] ),
    .B(\soc/cpu/timer[25] ),
    .C(\soc/cpu/timer[24] ),
    .D(\soc/cpu/timer[27] ),
    .Y(\soc/cpu/_01035_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05222_  (.A(\soc/cpu/_01032_ ),
    .B(\soc/cpu/_01033_ ),
    .C(\soc/cpu/_01034_ ),
    .D(\soc/cpu/_01035_ ),
    .Y(\soc/cpu/_01036_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05223_  (.A(\soc/cpu/_01031_ ),
    .B(\soc/cpu/_01036_ ),
    .Y(\soc/cpu/_01037_ ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_05224_  (.A(\soc/cpu/_01027_ ),
    .B(\soc/cpu/_01029_ ),
    .C(\soc/cpu/_01037_ ),
    .X(\soc/cpu/_01038_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05225_  (.A(\soc/cpu/_01023_ ),
    .B(\soc/cpu/_01025_ ),
    .C(\soc/cpu/_01026_ ),
    .D(\soc/cpu/_01038_ ),
    .Y(\soc/cpu/_01039_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05226_  (.A(\soc/cpu/timer[14] ),
    .B(\soc/cpu/_01005_ ),
    .Y(\soc/cpu/_01040_ ));
 sky130_fd_sc_hd__nor4b_2 \soc/cpu/_05227_  (.A(\soc/cpu/timer[16] ),
    .B(\soc/cpu/_01022_ ),
    .C(\soc/cpu/_01039_ ),
    .D_N(\soc/cpu/_01040_ ),
    .Y(\soc/cpu/_01041_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_05228_  (.A(\soc/cpu/_01019_ ),
    .B(\soc/cpu/_01021_ ),
    .C(\soc/cpu/_01041_ ),
    .X(\soc/cpu/_01042_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05229_  (.A(\soc/cpu/_01016_ ),
    .B(\soc/cpu/_01018_ ),
    .C(\soc/cpu/_01042_ ),
    .Y(\soc/cpu/_01043_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_05230_  (.A1(net876),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[0] ),
    .C1(_074_),
    .Y(\soc/cpu/_01044_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_05231_  (.A_N(net447),
    .B(\soc/cpu/_01043_ ),
    .C(\soc/cpu/_01044_ ),
    .Y(\soc/cpu/_00001_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05232_  (.A(\soc/cpu/mem_rdata_q[25] ),
    .B(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01045_ ));
 sky130_fd_sc_hd__o21bai_2 \soc/cpu/_05234_  (.A1(\soc/mem_rdata[25] ),
    .A2(net65),
    .B1_N(\soc/cpu/_01045_ ),
    .Y(\soc/cpu/_01047_ ));
 sky130_fd_sc_hd__inv_12 \soc/cpu/_05235_  (.A(\soc/cpu/mem_la_secondword ),
    .Y(\soc/cpu/_01048_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05237_  (.A(\soc/cpu/_01048_ ),
    .B(\soc/cpu/_00725_ ),
    .Y(\soc/cpu/_01050_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05238_  (.A0(\soc/cpu/mem_rdata_q[9] ),
    .A1(\soc/mem_rdata[9] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01051_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05240_  (.A1(\soc/cpu/_01047_ ),
    .A2(\soc/cpu/_01050_ ),
    .B1(\soc/cpu/_01051_ ),
    .B2(\soc/cpu/_01048_ ),
    .Y(\soc/cpu/_01053_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05241_  (.A(net65),
    .B(\soc/cpu/_01053_ ),
    .Y(\soc/cpu/_01054_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05242_  (.A(\soc/cpu/_01045_ ),
    .B(\soc/cpu/_01054_ ),
    .Y(\soc/cpu/_01055_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05243_  (.A(\soc/cpu/_01055_ ),
    .Y(\soc/cpu/_01056_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05244_  (.A(\soc/cpu/_00730_ ),
    .B(\soc/cpu/_00826_ ),
    .Y(\soc/cpu/_01057_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_05246_  (.A(\soc/cpu/mem_rdata_q[30] ),
    .B(\soc/cpu/_00721_ ),
    .X(\soc/cpu/_01059_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05247_  (.A1(\soc/mem_rdata[30] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01059_ ),
    .Y(\soc/cpu/_01060_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05248_  (.A0(\soc/cpu/mem_rdata_q[14] ),
    .A1(\soc/mem_rdata[14] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01061_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05249_  (.A1(net133),
    .A2(\soc/cpu/_01061_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01062_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05250_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01060_ ),
    .B1(\soc/cpu/_01062_ ),
    .Y(\soc/cpu/_01063_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_05251_  (.A1(\soc/cpu/mem_16bit_buffer[14] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01063_ ),
    .X(\soc/cpu/_01064_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05254_  (.A0(\soc/cpu/mem_rdata_q[13] ),
    .A1(\soc/mem_rdata[13] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01067_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_05255_  (.A(\soc/cpu/mem_rdata_q[29] ),
    .B(\soc/cpu/_00718_ ),
    .X(\soc/cpu/_01068_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05256_  (.A1(\soc/mem_rdata[29] ),
    .A2(\soc/cpu/_00721_ ),
    .B1(\soc/cpu/_01068_ ),
    .Y(\soc/cpu/_01069_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05257_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01069_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01070_ ));
 sky130_fd_sc_hd__o21bai_2 \soc/cpu/_05258_  (.A1(net133),
    .A2(\soc/cpu/_01067_ ),
    .B1_N(\soc/cpu/_01070_ ),
    .Y(\soc/cpu/_01071_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05259_  (.A1(\soc/cpu/mem_16bit_buffer[13] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01071_ ),
    .Y(\soc/cpu/_01072_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05260_  (.A0(\soc/mem_rdata[15] ),
    .A1(\soc/cpu/mem_rdata_q[15] ),
    .S(net65),
    .Y(\soc/cpu/_01073_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_05261_  (.A(\soc/cpu/mem_rdata_q[31] ),
    .B(net65),
    .X(\soc/cpu/_01074_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05262_  (.A1(\soc/mem_rdata[31] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01074_ ),
    .Y(\soc/cpu/_01075_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05263_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01075_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01076_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05264_  (.A1(net133),
    .A2(\soc/cpu/_01073_ ),
    .B1(\soc/cpu/_01076_ ),
    .Y(\soc/cpu/_01077_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_05265_  (.A1(\soc/cpu/mem_16bit_buffer[15] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01077_ ),
    .X(\soc/cpu/_01078_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05267_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01078_ ),
    .Y(\soc/cpu/_01080_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_05268_  (.A(\soc/cpu/_01064_ ),
    .B(\soc/cpu/_01080_ ),
    .Y(\soc/cpu/_01081_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05269_  (.A(\soc/cpu/mem_rdata_q[5] ),
    .B(net66),
    .Y(\soc/cpu/_01082_ ));
 sky130_fd_sc_hd__a21boi_2 \soc/cpu/_05270_  (.A1(\soc/mem_rdata[5] ),
    .A2(\soc/cpu/_00718_ ),
    .B1_N(\soc/cpu/_01082_ ),
    .Y(\soc/cpu/_01083_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05271_  (.A(\soc/cpu/mem_rdata_q[21] ),
    .B(net66),
    .X(\soc/cpu/_01084_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05272_  (.A1(\soc/mem_rdata[21] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01084_ ),
    .Y(\soc/cpu/_01085_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05273_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01085_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01086_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05274_  (.A1(net133),
    .A2(\soc/cpu/_01083_ ),
    .B1(\soc/cpu/_01086_ ),
    .Y(\soc/cpu/_01087_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05275_  (.A1(\soc/cpu/mem_16bit_buffer[5] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01087_ ),
    .Y(\soc/cpu/_01088_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05276_  (.A(\soc/cpu/mem_rdata_q[6] ),
    .B(net66),
    .Y(\soc/cpu/_01089_ ));
 sky130_fd_sc_hd__a21boi_2 \soc/cpu/_05277_  (.A1(\soc/mem_rdata[6] ),
    .A2(\soc/cpu/_00718_ ),
    .B1_N(\soc/cpu/_01089_ ),
    .Y(\soc/cpu/_01090_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05278_  (.A(\soc/cpu/mem_rdata_q[22] ),
    .B(net66),
    .X(\soc/cpu/_01091_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05279_  (.A1(\soc/mem_rdata[22] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01091_ ),
    .Y(\soc/cpu/_01092_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05280_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01092_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01093_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05281_  (.A1(net133),
    .A2(\soc/cpu/_01090_ ),
    .B1(\soc/cpu/_01093_ ),
    .Y(\soc/cpu/_01094_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05282_  (.A1(\soc/cpu/mem_16bit_buffer[6] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01094_ ),
    .Y(\soc/cpu/_01095_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05283_  (.A(\soc/cpu/mem_rdata_q[4] ),
    .B(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_01096_ ));
 sky130_fd_sc_hd__a21boi_2 \soc/cpu/_05284_  (.A1(\soc/mem_rdata[4] ),
    .A2(\soc/cpu/_00718_ ),
    .B1_N(\soc/cpu/_01096_ ),
    .Y(\soc/cpu/_01097_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05285_  (.A(\soc/cpu/_00713_ ),
    .B(\soc/cpu/_01097_ ),
    .Y(\soc/cpu/_01098_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05286_  (.A(\soc/cpu/mem_rdata_q[20] ),
    .B(net66),
    .X(\soc/cpu/_01099_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05287_  (.A1(\soc/mem_rdata[20] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01099_ ),
    .Y(\soc/cpu/_01100_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05288_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01100_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01101_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05289_  (.A1(\soc/cpu/mem_16bit_buffer[4] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01098_ ),
    .B2(\soc/cpu/_01101_ ),
    .Y(\soc/cpu/_01102_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05290_  (.A(\soc/cpu/_01088_ ),
    .B(\soc/cpu/_01095_ ),
    .C(\soc/cpu/_01102_ ),
    .Y(\soc/cpu/_01103_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05292_  (.A(\soc/mem_rdata[2] ),
    .B(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01105_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05293_  (.A(\soc/cpu/mem_rdata_q[2] ),
    .B(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_01106_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05294_  (.A1(\soc/cpu/_01105_ ),
    .A2(\soc/cpu/_01106_ ),
    .B1(\soc/cpu/_00713_ ),
    .Y(\soc/cpu/_01107_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05295_  (.A0(\soc/mem_rdata[18] ),
    .A1(\soc/cpu/mem_rdata_q[18] ),
    .S(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_01108_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05296_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01108_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01109_ ));
 sky130_fd_sc_hd__o22a_4 \soc/cpu/_05297_  (.A1(\soc/cpu/mem_16bit_buffer[2] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01107_ ),
    .B2(\soc/cpu/_01109_ ),
    .X(\soc/cpu/_01110_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05298_  (.A(\soc/cpu/mem_rdata_q[3] ),
    .B(net65),
    .Y(\soc/cpu/_01111_ ));
 sky130_fd_sc_hd__a21boi_2 \soc/cpu/_05299_  (.A1(\soc/mem_rdata[3] ),
    .A2(\soc/cpu/_00718_ ),
    .B1_N(\soc/cpu/_01111_ ),
    .Y(\soc/cpu/_01112_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05300_  (.A0(\soc/mem_rdata[19] ),
    .A1(\soc/cpu/mem_rdata_q[19] ),
    .S(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_01113_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05301_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01113_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01114_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05302_  (.A1(\soc/cpu/_00713_ ),
    .A2(\soc/cpu/_01112_ ),
    .B1(\soc/cpu/_01114_ ),
    .Y(\soc/cpu/_01115_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_05303_  (.A1(\soc/cpu/mem_16bit_buffer[3] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01115_ ),
    .X(\soc/cpu/_01116_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_05304_  (.A(\soc/cpu/_01103_ ),
    .B(\soc/cpu/_01110_ ),
    .C(\soc/cpu/_01116_ ),
    .Y(\soc/cpu/_01117_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05305_  (.A(\soc/cpu/_01081_ ),
    .B(\soc/cpu/_01117_ ),
    .Y(\soc/cpu/_01118_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05307_  (.A0(\soc/mem_rdata[12] ),
    .A1(\soc/cpu/mem_rdata_q[12] ),
    .S(\soc/cpu/_00721_ ),
    .Y(\soc/cpu/_01120_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05308_  (.A0(\soc/mem_rdata[28] ),
    .A1(\soc/cpu/mem_rdata_q[28] ),
    .S(net65),
    .Y(\soc/cpu/_01121_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05309_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01121_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01122_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05310_  (.A1(\soc/cpu/_00713_ ),
    .A2(\soc/cpu/_01120_ ),
    .B1(\soc/cpu/_01122_ ),
    .Y(\soc/cpu/_01123_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_05311_  (.A1(\soc/cpu/mem_16bit_buffer[12] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01123_ ),
    .X(\soc/cpu/_01124_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05312_  (.A0(\soc/cpu/mem_rdata_q[27] ),
    .A1(\soc/mem_rdata[27] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01125_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05313_  (.A(\soc/cpu/_00725_ ),
    .B(\soc/cpu/_01125_ ),
    .Y(\soc/cpu/_01126_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05314_  (.A(\soc/cpu/mem_rdata_q[11] ),
    .B(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01127_ ));
 sky130_fd_sc_hd__o21bai_2 \soc/cpu/_05315_  (.A1(\soc/mem_rdata[11] ),
    .A2(net66),
    .B1_N(\soc/cpu/_01127_ ),
    .Y(\soc/cpu/_01128_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05316_  (.A1(net133),
    .A2(\soc/cpu/_01128_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01129_ ));
 sky130_fd_sc_hd__o22a_4 \soc/cpu/_05317_  (.A1(\soc/cpu/mem_16bit_buffer[11] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01126_ ),
    .B2(\soc/cpu/_01129_ ),
    .X(\soc/cpu/_01130_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05318_  (.A(\soc/cpu/mem_rdata_q[8] ),
    .B(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01131_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_05319_  (.A1(\soc/mem_rdata[8] ),
    .A2(net65),
    .B1_N(\soc/cpu/_01131_ ),
    .Y(\soc/cpu/_01132_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05320_  (.A(net133),
    .B(\soc/cpu/_01132_ ),
    .Y(\soc/cpu/_01133_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05321_  (.A(\soc/cpu/mem_rdata_q[24] ),
    .B(net65),
    .X(\soc/cpu/_01134_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05322_  (.A1(\soc/mem_rdata[24] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01134_ ),
    .Y(\soc/cpu/_01135_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05323_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01135_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01136_ ));
 sky130_fd_sc_hd__o22a_4 \soc/cpu/_05324_  (.A1(\soc/cpu/mem_16bit_buffer[8] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01133_ ),
    .B2(\soc/cpu/_01136_ ),
    .X(\soc/cpu/_01137_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05325_  (.A(\soc/cpu/_00725_ ),
    .B(\soc/cpu/_01047_ ),
    .Y(\soc/cpu/_01138_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05326_  (.A1(net133),
    .A2(\soc/cpu/_01051_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01139_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05327_  (.A1(\soc/cpu/mem_16bit_buffer[9] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01138_ ),
    .B2(\soc/cpu/_01139_ ),
    .Y(\soc/cpu/_01140_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_05328_  (.A(\soc/cpu/mem_rdata_q[23] ),
    .B(net66),
    .X(\soc/cpu/_01141_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05329_  (.A1(\soc/mem_rdata[23] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01141_ ),
    .Y(\soc/cpu/_01142_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05330_  (.A0(\soc/cpu/mem_rdata_q[7] ),
    .A1(\soc/mem_rdata[7] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01143_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05331_  (.A1(net133),
    .A2(\soc/cpu/_01143_ ),
    .B1(\soc/cpu/_00716_ ),
    .X(\soc/cpu/_01144_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05332_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01142_ ),
    .B1(\soc/cpu/_01144_ ),
    .Y(\soc/cpu/_01145_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05333_  (.A1(\soc/cpu/mem_16bit_buffer[7] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01145_ ),
    .Y(\soc/cpu/_01146_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05334_  (.A0(\soc/cpu/mem_rdata_q[10] ),
    .A1(\soc/mem_rdata[10] ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01147_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05335_  (.A(net133),
    .B(\soc/cpu/_01147_ ),
    .Y(\soc/cpu/_01148_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05336_  (.A(\soc/cpu/mem_rdata_q[26] ),
    .B(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01149_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_05337_  (.A1(\soc/mem_rdata[26] ),
    .A2(net65),
    .B1_N(\soc/cpu/_01149_ ),
    .Y(\soc/cpu/_01150_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05338_  (.A1(\soc/cpu/_00725_ ),
    .A2(\soc/cpu/_01150_ ),
    .B1(\soc/cpu/_00716_ ),
    .Y(\soc/cpu/_01151_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05339_  (.A1(\soc/cpu/mem_16bit_buffer[10] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01148_ ),
    .B2(\soc/cpu/_01151_ ),
    .Y(\soc/cpu/_01152_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_05340_  (.A(\soc/cpu/_01140_ ),
    .B(\soc/cpu/_01146_ ),
    .C(\soc/cpu/_01152_ ),
    .X(\soc/cpu/_01153_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05341_  (.A_N(\soc/cpu/_01137_ ),
    .B(\soc/cpu/_01153_ ),
    .Y(\soc/cpu/_01154_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05342_  (.A(\soc/cpu/_01130_ ),
    .B(\soc/cpu/_01154_ ),
    .Y(\soc/cpu/_01155_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05343_  (.A(\soc/cpu/_01124_ ),
    .B(\soc/cpu/_01155_ ),
    .Y(\soc/cpu/_01156_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05345_  (.A1(\soc/cpu/_01118_ ),
    .A2(\soc/cpu/_01156_ ),
    .B1(\soc/cpu/_01072_ ),
    .Y(\soc/cpu/_01158_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_05346_  (.A(\soc/cpu/mem_do_prefetch ),
    .B(\soc/cpu/mem_do_rinst ),
    .Y(\soc/cpu/_01159_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_05347_  (.A(\soc/cpu/_01159_ ),
    .B(\soc/cpu/_00833_ ),
    .Y(\soc/cpu/_01160_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05348_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01160_ ),
    .Y(\soc/cpu/_01161_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05349_  (.A1(\soc/cpu/_01057_ ),
    .A2(\soc/cpu/_01158_ ),
    .B1(\soc/cpu/_01161_ ),
    .Y(\soc/cpu/_01162_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_05350_  (.A1(\soc/cpu/mem_16bit_buffer[13] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01071_ ),
    .X(\soc/cpu/_01163_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05351_  (.A1(\soc/cpu/mem_16bit_buffer[14] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01063_ ),
    .Y(\soc/cpu/_01164_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05352_  (.A(\soc/cpu/_01163_ ),
    .B(\soc/cpu/_01164_ ),
    .Y(\soc/cpu/_01165_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_05353_  (.A(\soc/cpu/_00825_ ),
    .B(\soc/cpu/_00737_ ),
    .Y(\soc/cpu/_01166_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05356_  (.A1(\soc/cpu/mem_16bit_buffer[15] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01077_ ),
    .Y(\soc/cpu/_01169_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_05357_  (.A(\soc/cpu/_01163_ ),
    .B(\soc/cpu/_01064_ ),
    .C(\soc/cpu/_01169_ ),
    .Y(\soc/cpu/_01170_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05358_  (.A1(\soc/cpu/mem_16bit_buffer[11] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01126_ ),
    .B2(\soc/cpu/_01129_ ),
    .Y(\soc/cpu/_01171_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05359_  (.A(\soc/cpu/_01171_ ),
    .B(\soc/cpu/_01153_ ),
    .X(\soc/cpu/_01172_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05360_  (.A(\soc/cpu/_01137_ ),
    .B(\soc/cpu/_01172_ ),
    .Y(\soc/cpu/_01173_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05361_  (.A(\soc/cpu/_01064_ ),
    .B(\soc/cpu/_01078_ ),
    .Y(\soc/cpu/_01174_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05362_  (.A1(\soc/cpu/_01170_ ),
    .A2(\soc/cpu/_01173_ ),
    .B1(\soc/cpu/_01174_ ),
    .Y(\soc/cpu/_01175_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05363_  (.A(\soc/cpu/_01110_ ),
    .B(\soc/cpu/_01175_ ),
    .Y(\soc/cpu/_01176_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05364_  (.A(\soc/cpu/_01081_ ),
    .B(\soc/cpu/_01124_ ),
    .Y(\soc/cpu/_01177_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05365_  (.A(\soc/cpu/_01171_ ),
    .B(\soc/cpu/_01177_ ),
    .Y(\soc/cpu/_01178_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05366_  (.A1(\soc/cpu/_01055_ ),
    .A2(\soc/cpu/_01152_ ),
    .B1(\soc/cpu/_01178_ ),
    .Y(\soc/cpu/_01179_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_05367_  (.A1(\soc/cpu/_01137_ ),
    .A2(\soc/cpu/_01172_ ),
    .B1(\soc/cpu/_01170_ ),
    .Y(\soc/cpu/_01180_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05368_  (.A(\soc/cpu/_01124_ ),
    .B(\soc/cpu/_01180_ ),
    .Y(\soc/cpu/_01181_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_05370_  (.A(\soc/cpu/_01163_ ),
    .B(\soc/cpu/_01078_ ),
    .Y(\soc/cpu/_01183_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05372_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01064_ ),
    .Y(\soc/cpu/_01185_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05373_  (.A1(\soc/cpu/_01124_ ),
    .A2(\soc/cpu/_01183_ ),
    .B1(\soc/cpu/_01185_ ),
    .Y(\soc/cpu/_01186_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05374_  (.A(\soc/cpu/_01176_ ),
    .B(\soc/cpu/_01179_ ),
    .C(\soc/cpu/_01181_ ),
    .D(\soc/cpu/_01186_ ),
    .Y(\soc/cpu/_01187_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_05375_  (.A1(\soc/cpu/_01055_ ),
    .A2(\soc/cpu/_01165_ ),
    .B1(\soc/cpu/_01166_ ),
    .C1(\soc/cpu/_01187_ ),
    .Y(\soc/cpu/_01188_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05376_  (.A(\soc/cpu/_00825_ ),
    .B(\soc/cpu/_00737_ ),
    .Y(\soc/cpu/_01189_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05378_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01064_ ),
    .Y(\soc/cpu/_01191_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05379_  (.A(\soc/cpu/_01189_ ),
    .B(\soc/cpu/_01191_ ),
    .Y(\soc/cpu/_01192_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05380_  (.A(\soc/cpu/_00825_ ),
    .B(\soc/cpu/_00826_ ),
    .Y(\soc/cpu/_01193_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05381_  (.A(\soc/cpu/_01163_ ),
    .B(\soc/cpu/_01164_ ),
    .Y(\soc/cpu/_01194_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05382_  (.A(\soc/cpu/_01183_ ),
    .B(\soc/cpu/_01194_ ),
    .Y(\soc/cpu/_01195_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05383_  (.A(\soc/cpu/_01193_ ),
    .B(\soc/cpu/_01195_ ),
    .Y(\soc/cpu/_01196_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05384_  (.A1(\soc/cpu/_01192_ ),
    .A2(\soc/cpu/_01196_ ),
    .B1(\soc/cpu/_01124_ ),
    .Y(\soc/cpu/_01197_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_05385_  (.A(\soc/cpu/_00730_ ),
    .B(\soc/cpu/_00737_ ),
    .Y(\soc/cpu/_01198_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05386_  (.A(\soc/cpu/_01055_ ),
    .B(\soc/cpu/_01198_ ),
    .C(\soc/cpu/_01195_ ),
    .Y(\soc/cpu/_01199_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_05387_  (.A(\soc/cpu/_01188_ ),
    .B(\soc/cpu/_01197_ ),
    .C(\soc/cpu/_01199_ ),
    .X(\soc/cpu/_01200_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05388_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_00963_ ),
    .Y(\soc/cpu/_01201_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_05390_  (.A1(\soc/cpu/_01056_ ),
    .A2(\soc/cpu/_01162_ ),
    .B1(\soc/cpu/_01200_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00051_ ));
 sky130_fd_sc_hd__o22a_2 \soc/cpu/_05393_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01147_ ),
    .B1(\soc/cpu/_01150_ ),
    .B2(\soc/cpu/_01050_ ),
    .X(\soc/cpu/_01205_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05394_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01205_ ),
    .B1(\soc/cpu/_01149_ ),
    .Y(\soc/cpu/_01206_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05395_  (.A(\soc/cpu/_01206_ ),
    .Y(\soc/cpu/_01207_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05396_  (.A(\soc/cpu/_01110_ ),
    .B(\soc/cpu/_01183_ ),
    .Y(\soc/cpu/_01208_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05397_  (.A1(\soc/cpu/_01169_ ),
    .A2(\soc/cpu/_01146_ ),
    .B1(\soc/cpu/_01208_ ),
    .Y(\soc/cpu/_01209_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/_05398_  (.A1(\soc/cpu/mem_16bit_buffer[5] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01087_ ),
    .X(\soc/cpu/_01210_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05399_  (.A(\soc/cpu/_01164_ ),
    .B(\soc/cpu/_01183_ ),
    .Y(\soc/cpu/_01211_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/_05400_  (.A1(\soc/cpu/mem_16bit_buffer[7] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01145_ ),
    .X(\soc/cpu/_01212_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/_05401_  (.A1(\soc/cpu/_01210_ ),
    .A2(\soc/cpu/_01191_ ),
    .B1(\soc/cpu/_01211_ ),
    .B2(\soc/cpu/_01212_ ),
    .C1(\soc/cpu/_01198_ ),
    .Y(\soc/cpu/_01213_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05402_  (.A1(\soc/cpu/_01195_ ),
    .A2(\soc/cpu/_01207_ ),
    .B1(\soc/cpu/_01213_ ),
    .Y(\soc/cpu/_01214_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05403_  (.A1(\soc/cpu/mem_16bit_buffer[12] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01123_ ),
    .Y(\soc/cpu/_01215_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05405_  (.A(\soc/cpu/_01215_ ),
    .B(\soc/cpu/_01170_ ),
    .Y(\soc/cpu/_01217_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05406_  (.A(\soc/cpu/_01088_ ),
    .B(\soc/cpu/_01181_ ),
    .Y(\soc/cpu/_01218_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05407_  (.A1(\soc/cpu/_01175_ ),
    .A2(\soc/cpu/_01217_ ),
    .B1(\soc/cpu/_01218_ ),
    .Y(\soc/cpu/_01219_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05408_  (.A1(\soc/cpu/_01152_ ),
    .A2(\soc/cpu/_01206_ ),
    .B1(\soc/cpu/_01178_ ),
    .Y(\soc/cpu/_01220_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05409_  (.A1(\soc/cpu/_01165_ ),
    .A2(\soc/cpu/_01206_ ),
    .B1(\soc/cpu/_01166_ ),
    .Y(\soc/cpu/_01221_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05410_  (.A1(\soc/cpu/_01186_ ),
    .A2(\soc/cpu/_01219_ ),
    .A3(\soc/cpu/_01220_ ),
    .B1(\soc/cpu/_01221_ ),
    .Y(\soc/cpu/_01222_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05411_  (.A1(\soc/cpu/_01192_ ),
    .A2(\soc/cpu/_01209_ ),
    .B1(\soc/cpu/_01214_ ),
    .C1(\soc/cpu/_01222_ ),
    .Y(\soc/cpu/_01223_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_05412_  (.A1(\soc/cpu/_01162_ ),
    .A2(\soc/cpu/_01207_ ),
    .B1(\soc/cpu/_01223_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00052_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05413_  (.A1(\soc/cpu/_01050_ ),
    .A2(\soc/cpu/_01125_ ),
    .B1(\soc/cpu/_01128_ ),
    .B2(\soc/cpu/_01048_ ),
    .Y(\soc/cpu/_01224_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05414_  (.A0(\soc/cpu/mem_rdata_q[27] ),
    .A1(\soc/cpu/_01224_ ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01225_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05415_  (.A(\soc/cpu/_01170_ ),
    .B(\soc/cpu/_01173_ ),
    .Y(\soc/cpu/_01226_ ));
 sky130_fd_sc_hd__o22a_4 \soc/cpu/_05417_  (.A1(\soc/cpu/mem_16bit_buffer[10] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01148_ ),
    .B2(\soc/cpu/_01151_ ),
    .X(\soc/cpu/_01228_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05418_  (.A(\soc/cpu/_01228_ ),
    .B(\soc/cpu/_01225_ ),
    .Y(\soc/cpu/_01229_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05419_  (.A(\soc/cpu/_01178_ ),
    .B(\soc/cpu/_01229_ ),
    .Y(\soc/cpu/_01230_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_05420_  (.A1(\soc/cpu/_01095_ ),
    .A2(\soc/cpu/_01174_ ),
    .B1(\soc/cpu/_01181_ ),
    .C1(\soc/cpu/_01186_ ),
    .D1(\soc/cpu/_01230_ ),
    .Y(\soc/cpu/_01231_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05421_  (.A1(\soc/cpu/_01116_ ),
    .A2(\soc/cpu/_01226_ ),
    .B1(\soc/cpu/_01231_ ),
    .Y(\soc/cpu/_01232_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_05422_  (.A(\soc/cpu/_00730_ ),
    .B(\soc/cpu/_00826_ ),
    .Y(\soc/cpu/_01233_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05423_  (.A1(\soc/cpu/_01185_ ),
    .A2(\soc/cpu/_01225_ ),
    .B1(\soc/cpu/_01232_ ),
    .C1(\soc/cpu/_01233_ ),
    .Y(\soc/cpu/_01234_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05424_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01169_ ),
    .Y(\soc/cpu/_01235_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05425_  (.A(\soc/cpu/_01064_ ),
    .B(\soc/cpu/_01235_ ),
    .Y(\soc/cpu/_01236_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05426_  (.A(\soc/cpu/_01198_ ),
    .B(\soc/cpu/_01236_ ),
    .Y(\soc/cpu/_01237_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05427_  (.A(\soc/cpu/_01078_ ),
    .B(\soc/cpu/_01192_ ),
    .Y(\soc/cpu/_01238_ ));
 sky130_fd_sc_hd__a21boi_0 \soc/cpu/_05428_  (.A1(\soc/cpu/_01237_ ),
    .A2(\soc/cpu/_01238_ ),
    .B1_N(\soc/cpu/_01137_ ),
    .Y(\soc/cpu/_01239_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05429_  (.A(\soc/cpu/_01198_ ),
    .B(\soc/cpu/_01195_ ),
    .Y(\soc/cpu/_01240_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05430_  (.A1(\soc/cpu/mem_16bit_buffer[3] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01115_ ),
    .Y(\soc/cpu/_01241_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05431_  (.A(\soc/cpu/_01241_ ),
    .B(\soc/cpu/_01235_ ),
    .Y(\soc/cpu/_01242_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05432_  (.A(\soc/cpu/_01192_ ),
    .B(\soc/cpu/_01242_ ),
    .Y(\soc/cpu/_01243_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05433_  (.A1(\soc/cpu/_01225_ ),
    .A2(\soc/cpu/_01240_ ),
    .B1(\soc/cpu/_01243_ ),
    .Y(\soc/cpu/_01244_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05434_  (.A(\soc/cpu/_01234_ ),
    .B(\soc/cpu/_01239_ ),
    .C(\soc/cpu/_01244_ ),
    .Y(\soc/cpu/_01245_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05435_  (.A1(\soc/cpu/_01162_ ),
    .A2(\soc/cpu/_01225_ ),
    .B1(\soc/cpu/_01245_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00053_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05436_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01120_ ),
    .B1(\soc/cpu/_01121_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01246_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05437_  (.A0(\soc/cpu/mem_rdata_q[28] ),
    .A1(\soc/cpu/_01246_ ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01247_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05438_  (.A(\soc/cpu/_01185_ ),
    .B(\soc/cpu/_01166_ ),
    .Y(\soc/cpu/_01248_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_05439_  (.A(\soc/cpu/_01162_ ),
    .B(\soc/cpu/_01248_ ),
    .X(\soc/cpu/_01249_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_05440_  (.A(\soc/cpu/_01102_ ),
    .B(\soc/cpu/_01170_ ),
    .C(\soc/cpu/_01173_ ),
    .X(\soc/cpu/_01250_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05441_  (.A(\soc/cpu/_01228_ ),
    .B(\soc/cpu/_01247_ ),
    .Y(\soc/cpu/_01251_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05442_  (.A1(\soc/cpu/_01174_ ),
    .A2(\soc/cpu/_01235_ ),
    .B1(\soc/cpu/_01215_ ),
    .Y(\soc/cpu/_01252_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05443_  (.A1(\soc/cpu/_01178_ ),
    .A2(\soc/cpu/_01251_ ),
    .B1(\soc/cpu/_01252_ ),
    .Y(\soc/cpu/_01253_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05444_  (.A(\soc/cpu/_01165_ ),
    .B(\soc/cpu/_01166_ ),
    .Y(\soc/cpu/_01254_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05445_  (.A1(\soc/cpu/_01181_ ),
    .A2(\soc/cpu/_01250_ ),
    .A3(\soc/cpu/_01253_ ),
    .B1(\soc/cpu/_01254_ ),
    .Y(\soc/cpu/_01255_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05446_  (.A1(\soc/cpu/_01140_ ),
    .A2(\soc/cpu/_01237_ ),
    .B1(\soc/cpu/_01240_ ),
    .B2(\soc/cpu/_01247_ ),
    .Y(\soc/cpu/_01256_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05447_  (.A1(\soc/cpu/_01255_ ),
    .A2(\soc/cpu/_01256_ ),
    .B1(\soc/cpu/_01160_ ),
    .Y(\soc/cpu/_01257_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05448_  (.A1(\soc/cpu/_01247_ ),
    .A2(\soc/cpu/_01249_ ),
    .B1(\soc/cpu/_01257_ ),
    .Y(\soc/cpu/_00054_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05449_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01067_ ),
    .B1(\soc/cpu/_01069_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01258_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05450_  (.A1(\soc/cpu/_00721_ ),
    .A2(\soc/cpu/_01258_ ),
    .B1(\soc/cpu/_01068_ ),
    .Y(\soc/cpu/_01259_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05451_  (.A(\soc/cpu/_01185_ ),
    .B(\soc/cpu/_01233_ ),
    .Y(\soc/cpu/_01260_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05452_  (.A(\soc/cpu/_01260_ ),
    .B(\soc/cpu/_01178_ ),
    .Y(\soc/cpu/_01261_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05453_  (.A1(\soc/cpu/_01240_ ),
    .A2(\soc/cpu/_01261_ ),
    .B1(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_01262_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_05454_  (.A(\soc/cpu/_01249_ ),
    .SLEEP(\soc/cpu/_01262_ ),
    .X(\soc/cpu/_01263_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05455_  (.A1(\soc/cpu/_01064_ ),
    .A2(\soc/cpu/_01183_ ),
    .B1(\soc/cpu/_01124_ ),
    .Y(\soc/cpu/_01264_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05456_  (.A(\soc/cpu/_01254_ ),
    .B(\soc/cpu/_01264_ ),
    .Y(\soc/cpu/_01265_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05457_  (.A1(\soc/cpu/_01152_ ),
    .A2(\soc/cpu/_01260_ ),
    .A3(\soc/cpu/_01178_ ),
    .B1(\soc/cpu/_01265_ ),
    .Y(\soc/cpu/_01266_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05458_  (.A1(\soc/cpu/_01152_ ),
    .A2(\soc/cpu/_01237_ ),
    .B1(\soc/cpu/_01266_ ),
    .Y(\soc/cpu/_01267_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05459_  (.A(\soc/cpu/_01160_ ),
    .B(\soc/cpu/_01267_ ),
    .Y(\soc/cpu/_01268_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05460_  (.A1(\soc/cpu/_01259_ ),
    .A2(\soc/cpu/_01263_ ),
    .B1(\soc/cpu/_01268_ ),
    .Y(\soc/cpu/_00055_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05462_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01061_ ),
    .B1(\soc/cpu/_01060_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01270_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05463_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01270_ ),
    .B1(\soc/cpu/_01059_ ),
    .Y(\soc/cpu/_01271_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05464_  (.A(\soc/cpu/_01130_ ),
    .B(\soc/cpu/_01228_ ),
    .Y(\soc/cpu/_01272_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05465_  (.A(\soc/cpu/_01124_ ),
    .B(\soc/cpu/_01272_ ),
    .Y(\soc/cpu/_01273_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05466_  (.A(\soc/cpu/_01088_ ),
    .B(\soc/cpu/_01095_ ),
    .C(\soc/cpu/_01273_ ),
    .Y(\soc/cpu/_01274_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05467_  (.A1(\soc/cpu/_01215_ ),
    .A2(\soc/cpu/_01171_ ),
    .B1(\soc/cpu/_01152_ ),
    .Y(\soc/cpu/_01275_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05468_  (.A(\soc/cpu/_01272_ ),
    .B(\soc/cpu/_01275_ ),
    .Y(\soc/cpu/_01276_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05469_  (.A(\soc/cpu/_01274_ ),
    .B(\soc/cpu/_01276_ ),
    .Y(\soc/cpu/_01277_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05470_  (.A1(\soc/cpu/_01081_ ),
    .A2(\soc/cpu/_01166_ ),
    .A3(\soc/cpu/_01277_ ),
    .B1(\soc/cpu/_01265_ ),
    .Y(\soc/cpu/_01278_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05471_  (.A1(\soc/cpu/_01263_ ),
    .A2(\soc/cpu/_01271_ ),
    .B1(\soc/cpu/_01278_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00056_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_05472_  (.A(\soc/cpu/_01233_ ),
    .B(\soc/cpu/_01174_ ),
    .Y(\soc/cpu/_01279_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05473_  (.A(\soc/cpu/_01078_ ),
    .B(\soc/cpu/_01194_ ),
    .Y(\soc/cpu/_01280_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05474_  (.A(\soc/cpu/_00730_ ),
    .B(\soc/cpu/_01280_ ),
    .Y(\soc/cpu/_01281_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05475_  (.A(\soc/cpu/_01279_ ),
    .B(\soc/cpu/_01281_ ),
    .Y(\soc/cpu/_01282_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05476_  (.A(\soc/cpu/_01201_ ),
    .B(\soc/cpu/_01282_ ),
    .Y(\soc/cpu/_01283_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05478_  (.A(net65),
    .B(\soc/cpu/_01137_ ),
    .Y(\soc/cpu/_01285_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05479_  (.A(\soc/cpu/_01160_ ),
    .B(\soc/cpu/_01279_ ),
    .Y(\soc/cpu/_01286_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_05480_  (.A1(\soc/cpu/_01131_ ),
    .A2(\soc/cpu/_01283_ ),
    .A3(\soc/cpu/_01285_ ),
    .B1(\soc/cpu/_01286_ ),
    .B2(\soc/cpu/_01241_ ),
    .Y(\soc/cpu/_00059_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05481_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_01140_ ),
    .Y(\soc/cpu/_01287_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05482_  (.A1(\soc/cpu/mem_rdata_q[9] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01287_ ),
    .Y(\soc/cpu/_01288_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/_05483_  (.A1(\soc/cpu/mem_16bit_buffer[6] ),
    .A2(\soc/cpu/_00716_ ),
    .B1(\soc/cpu/_01094_ ),
    .X(\soc/cpu/_01289_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05484_  (.A(\soc/cpu/_01193_ ),
    .B(\soc/cpu/_01280_ ),
    .Y(\soc/cpu/_01290_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05485_  (.A(\soc/cpu/_01279_ ),
    .Y(\soc/cpu/_01291_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_05487_  (.A1(\soc/cpu/_01189_ ),
    .A2(\soc/cpu/_01140_ ),
    .A3(\soc/cpu/_01280_ ),
    .B1(\soc/cpu/_01291_ ),
    .B2(\soc/cpu/_01102_ ),
    .Y(\soc/cpu/_01293_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05488_  (.A1(\soc/cpu/_01289_ ),
    .A2(\soc/cpu/_01290_ ),
    .B1(\soc/cpu/_01293_ ),
    .Y(\soc/cpu/_01294_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05489_  (.A1(\soc/cpu/_01283_ ),
    .A2(\soc/cpu/_01288_ ),
    .B1(\soc/cpu/_01294_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00060_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05490_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_01152_ ),
    .Y(\soc/cpu/_01295_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05491_  (.A1(\soc/cpu/mem_rdata_q[10] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01295_ ),
    .Y(\soc/cpu/_01296_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05492_  (.A(\soc/cpu/_01228_ ),
    .B(\soc/cpu/_01283_ ),
    .Y(\soc/cpu/_01297_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05493_  (.A1(\soc/cpu/_01283_ ),
    .A2(\soc/cpu/_01296_ ),
    .B1(\soc/cpu/_01297_ ),
    .Y(\soc/cpu/_00036_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05494_  (.A1(\soc/cpu/_00826_ ),
    .A2(\soc/cpu/_01174_ ),
    .B1(\soc/cpu/_00825_ ),
    .Y(\soc/cpu/_01298_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05496_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01130_ ),
    .Y(\soc/cpu/_01300_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_05497_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01281_ ),
    .A3(\soc/cpu/_01298_ ),
    .B1(\soc/cpu/_01300_ ),
    .Y(\soc/cpu/_01301_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05499_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_01303_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05500_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01171_ ),
    .B1(\soc/cpu/_01303_ ),
    .Y(\soc/cpu/_01304_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05501_  (.A1(\soc/cpu/_01160_ ),
    .A2(\soc/cpu/_01301_ ),
    .B1(\soc/cpu/_01304_ ),
    .Y(\soc/cpu/_01305_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05502_  (.A(\soc/cpu/_01130_ ),
    .B(\soc/cpu/_01283_ ),
    .Y(\soc/cpu/_01306_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05503_  (.A1(\soc/cpu/_01127_ ),
    .A2(\soc/cpu/_01305_ ),
    .B1(\soc/cpu/_01306_ ),
    .Y(\soc/cpu/_00037_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05505_  (.A(net66),
    .B(\soc/cpu/_01215_ ),
    .Y(\soc/cpu/_01308_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05506_  (.A1(\soc/cpu/mem_rdata_q[12] ),
    .A2(net66),
    .B1(\soc/cpu/_01308_ ),
    .Y(\soc/cpu/_01309_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05507_  (.A(\soc/cpu/_01215_ ),
    .B(\soc/cpu/_01272_ ),
    .Y(\soc/cpu/_01310_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05508_  (.A1(\soc/cpu/_01088_ ),
    .A2(\soc/cpu/_01095_ ),
    .B1(\soc/cpu/_01273_ ),
    .Y(\soc/cpu/_01311_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05509_  (.A(\soc/cpu/_01081_ ),
    .B(\soc/cpu/_01311_ ),
    .Y(\soc/cpu/_01312_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05510_  (.A1(\soc/cpu/_01309_ ),
    .A2(\soc/cpu/_01310_ ),
    .B1(\soc/cpu/_01312_ ),
    .Y(\soc/cpu/_01313_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05511_  (.A1(\soc/cpu/_01110_ ),
    .A2(\soc/cpu/_01180_ ),
    .B1(\soc/cpu/_01313_ ),
    .Y(\soc/cpu/_01314_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05512_  (.A1(\soc/cpu/_01072_ ),
    .A2(\soc/cpu/_01174_ ),
    .B1(\soc/cpu/_01314_ ),
    .Y(\soc/cpu/_01315_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05513_  (.A1(\soc/cpu/_01189_ ),
    .A2(\soc/cpu/_01211_ ),
    .B1(\soc/cpu/_01240_ ),
    .B2(\soc/cpu/_01309_ ),
    .Y(\soc/cpu/_01316_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05514_  (.A1(\soc/cpu/_01260_ ),
    .A2(\soc/cpu/_01315_ ),
    .B1(\soc/cpu/_01316_ ),
    .Y(\soc/cpu/_01317_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05515_  (.A1(\soc/cpu/_01249_ ),
    .A2(\soc/cpu/_01309_ ),
    .B1(\soc/cpu/_01317_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00038_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05516_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_01072_ ),
    .Y(\soc/cpu/_01318_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05517_  (.A1(\soc/cpu/mem_rdata_q[13] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01318_ ),
    .Y(\soc/cpu/_01319_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05518_  (.A(\soc/cpu/_01124_ ),
    .B(\soc/cpu/_01228_ ),
    .C(\soc/cpu/_01319_ ),
    .Y(\soc/cpu/_01320_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05519_  (.A(\soc/cpu/_01081_ ),
    .B(\soc/cpu/_01130_ ),
    .C(\soc/cpu/_01320_ ),
    .Y(\soc/cpu/_01321_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05520_  (.A1(\soc/cpu/_01095_ ),
    .A2(\soc/cpu/_01273_ ),
    .B1(\soc/cpu/_01321_ ),
    .Y(\soc/cpu/_01322_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05521_  (.A1(\soc/cpu/_01116_ ),
    .A2(\soc/cpu/_01180_ ),
    .B1(\soc/cpu/_01322_ ),
    .Y(\soc/cpu/_01323_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05522_  (.A(\soc/cpu/_01254_ ),
    .B(\soc/cpu/_01323_ ),
    .Y(\soc/cpu/_01324_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05523_  (.A1(\soc/cpu/_01195_ ),
    .A2(\soc/cpu/_01319_ ),
    .B1(\soc/cpu/_01236_ ),
    .C1(\soc/cpu/_01193_ ),
    .Y(\soc/cpu/_01325_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05524_  (.A(\soc/cpu/_01192_ ),
    .B(\soc/cpu/_01324_ ),
    .C(\soc/cpu/_01325_ ),
    .Y(\soc/cpu/_01326_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05525_  (.A1(\soc/cpu/_01249_ ),
    .A2(\soc/cpu/_01319_ ),
    .B1(\soc/cpu/_01326_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00039_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05526_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01164_ ),
    .C(\soc/cpu/_01078_ ),
    .Y(\soc/cpu/_01327_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05527_  (.A(\soc/cpu/_01327_ ),
    .B(\soc/cpu/_01173_ ),
    .Y(\soc/cpu/_01328_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05528_  (.A(\soc/cpu/_01081_ ),
    .B(\soc/cpu/_01274_ ),
    .Y(\soc/cpu/_01329_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05529_  (.A1(\soc/cpu/_01102_ ),
    .A2(\soc/cpu/_01328_ ),
    .B1(\soc/cpu/_01310_ ),
    .B2(\soc/cpu/_01329_ ),
    .Y(\soc/cpu/_01330_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05530_  (.A(\soc/cpu/_01057_ ),
    .B(\soc/cpu/_01158_ ),
    .Y(\soc/cpu/_01331_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05532_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_01164_ ),
    .Y(\soc/cpu/_01333_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05533_  (.A1(\soc/cpu/mem_rdata_q[14] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01333_ ),
    .Y(\soc/cpu/_01334_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05534_  (.A1(\soc/cpu/_01331_ ),
    .A2(\soc/cpu/_01240_ ),
    .B1(\soc/cpu/_01334_ ),
    .Y(\soc/cpu/_01335_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05535_  (.A1(\soc/cpu/_01260_ ),
    .A2(\soc/cpu/_01330_ ),
    .B1(\soc/cpu/_01335_ ),
    .Y(\soc/cpu/_01336_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05536_  (.A1(\soc/cpu/_01165_ ),
    .A2(\soc/cpu/_01329_ ),
    .B1(\soc/cpu/_01233_ ),
    .Y(\soc/cpu/_01337_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05537_  (.A(\soc/cpu/_01161_ ),
    .B(\soc/cpu/_01337_ ),
    .Y(\soc/cpu/_01338_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05538_  (.A1(\soc/cpu/_01201_ ),
    .A2(\soc/cpu/_01336_ ),
    .B1(\soc/cpu/_01338_ ),
    .B2(\soc/cpu/_01334_ ),
    .Y(\soc/cpu/_00040_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_05539_  (.A(\soc/cpu/_01201_ ),
    .B(\soc/cpu/_01233_ ),
    .C(\soc/cpu/_01328_ ),
    .Y(\soc/cpu/_01339_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05540_  (.A(net66),
    .B(\soc/cpu/_01169_ ),
    .Y(\soc/cpu/_01340_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05541_  (.A1(\soc/cpu/mem_rdata_q[15] ),
    .A2(net66),
    .B1(\soc/cpu/_01339_ ),
    .C1(\soc/cpu/_01340_ ),
    .Y(\soc/cpu/_01341_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05542_  (.A1(\soc/cpu/_01088_ ),
    .A2(\soc/cpu/_01339_ ),
    .B1(\soc/cpu/_01341_ ),
    .Y(\soc/cpu/_00041_ ));
 sky130_fd_sc_hd__o22a_2 \soc/cpu/_05543_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_00724_ ),
    .B1(\soc/cpu/_00727_ ),
    .B2(\soc/cpu/_01050_ ),
    .X(\soc/cpu/_01342_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05544_  (.A(net66),
    .B(\soc/cpu/_01342_ ),
    .Y(\soc/cpu/_01343_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05545_  (.A1(\soc/cpu/mem_rdata_q[16] ),
    .A2(net66),
    .B1(\soc/cpu/_01339_ ),
    .C1(\soc/cpu/_01343_ ),
    .Y(\soc/cpu/_01344_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05546_  (.A1(\soc/cpu/_01095_ ),
    .A2(\soc/cpu/_01339_ ),
    .B1(\soc/cpu/_01344_ ),
    .Y(\soc/cpu/_00042_ ));
 sky130_fd_sc_hd__o22a_2 \soc/cpu/_05547_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_00733_ ),
    .B1(\soc/cpu/_00734_ ),
    .B2(\soc/cpu/_01050_ ),
    .X(\soc/cpu/_01345_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05548_  (.A(net66),
    .B(\soc/cpu/_01345_ ),
    .Y(\soc/cpu/_01346_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05549_  (.A1(\soc/cpu/mem_rdata_q[17] ),
    .A2(net66),
    .B1(\soc/cpu/_01346_ ),
    .Y(\soc/cpu/_01347_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05550_  (.A(\soc/cpu/_01124_ ),
    .B(\soc/cpu/_01339_ ),
    .Y(\soc/cpu/_01348_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05551_  (.A1(\soc/cpu/_01339_ ),
    .A2(\soc/cpu/_01347_ ),
    .B1(\soc/cpu/_01348_ ),
    .Y(\soc/cpu/_00043_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05552_  (.A(\soc/cpu/_01105_ ),
    .B(\soc/cpu/_01106_ ),
    .Y(\soc/cpu/_01349_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05553_  (.A(\soc/cpu/_01050_ ),
    .B(\soc/cpu/_01108_ ),
    .Y(\soc/cpu/_01350_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_05554_  (.A1(\soc/cpu/mem_la_secondword ),
    .A2(\soc/cpu/_01349_ ),
    .B1(\soc/cpu/_01350_ ),
    .Y(\soc/cpu/_01351_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05555_  (.A(net66),
    .B(\soc/cpu/_01351_ ),
    .Y(\soc/cpu/_01352_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05556_  (.A1(\soc/cpu/mem_rdata_q[18] ),
    .A2(net66),
    .B1(\soc/cpu/_01352_ ),
    .Y(\soc/cpu/_01353_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05557_  (.A1(\soc/cpu/_01339_ ),
    .A2(\soc/cpu/_01353_ ),
    .B1(\soc/cpu/_01348_ ),
    .Y(\soc/cpu/_00044_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05558_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01112_ ),
    .B1(\soc/cpu/_01113_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01354_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05559_  (.A0(\soc/cpu/mem_rdata_q[19] ),
    .A1(\soc/cpu/_01354_ ),
    .S(\soc/cpu/_00718_ ),
    .Y(\soc/cpu/_01355_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05560_  (.A1(\soc/cpu/_01339_ ),
    .A2(\soc/cpu/_01355_ ),
    .B1(\soc/cpu/_01348_ ),
    .Y(\soc/cpu/_00045_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05561_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01097_ ),
    .B1(\soc/cpu/_01100_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01356_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05562_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01356_ ),
    .B1(\soc/cpu/_01099_ ),
    .Y(\soc/cpu/_01357_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05563_  (.A(\soc/cpu/_01164_ ),
    .B(\soc/cpu/_01235_ ),
    .Y(\soc/cpu/_01358_ ));
 sky130_fd_sc_hd__a311oi_2 \soc/cpu/_05564_  (.A1(\soc/cpu/_01081_ ),
    .A2(\soc/cpu/_01117_ ),
    .A3(\soc/cpu/_01156_ ),
    .B1(\soc/cpu/_01358_ ),
    .C1(\soc/cpu/_01189_ ),
    .Y(\soc/cpu/_01359_ ));
 sky130_fd_sc_hd__a2111oi_2 \soc/cpu/_05565_  (.A1(\soc/cpu/_01185_ ),
    .A2(\soc/cpu/_01166_ ),
    .B1(\soc/cpu/_01279_ ),
    .C1(\soc/cpu/_01359_ ),
    .D1(\soc/cpu/_01161_ ),
    .Y(\soc/cpu/_01360_ ));
 sky130_fd_sc_hd__a21boi_1 \soc/cpu/_05566_  (.A1(\soc/cpu/_01235_ ),
    .A2(\soc/cpu/_01198_ ),
    .B1_N(\soc/cpu/_01360_ ),
    .Y(\soc/cpu/_01361_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05567_  (.A(\soc/cpu/_01130_ ),
    .B(\soc/cpu/_01152_ ),
    .Y(\soc/cpu/_01362_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_05568_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01164_ ),
    .C(\soc/cpu/_01078_ ),
    .Y(\soc/cpu/_01363_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05569_  (.A1(\soc/cpu/_01362_ ),
    .A2(\soc/cpu/_01357_ ),
    .B1(\soc/cpu/_01363_ ),
    .Y(\soc/cpu/_01364_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05570_  (.A1(\soc/cpu/_01110_ ),
    .A2(\soc/cpu/_01362_ ),
    .B1(\soc/cpu/_01364_ ),
    .Y(\soc/cpu/_01365_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05571_  (.A(\soc/cpu/_01181_ ),
    .B(\soc/cpu/_01208_ ),
    .C(\soc/cpu/_01365_ ),
    .Y(\soc/cpu/_01366_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05572_  (.A1(\soc/cpu/_01064_ ),
    .A2(\soc/cpu/_01078_ ),
    .B1(\soc/cpu/_01254_ ),
    .Y(\soc/cpu/_01367_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05573_  (.A(\soc/cpu/_01160_ ),
    .B(\soc/cpu/_01366_ ),
    .C(\soc/cpu/_01367_ ),
    .Y(\soc/cpu/_01368_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05574_  (.A1(\soc/cpu/_01357_ ),
    .A2(\soc/cpu/_01361_ ),
    .B1(\soc/cpu/_01368_ ),
    .Y(\soc/cpu/_00046_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05575_  (.A1(\soc/cpu/_01050_ ),
    .A2(\soc/cpu/_01085_ ),
    .B1(\soc/cpu/_01083_ ),
    .B2(\soc/cpu/_01048_ ),
    .Y(\soc/cpu/_01369_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05576_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01369_ ),
    .B1(\soc/cpu/_01084_ ),
    .Y(\soc/cpu/_01370_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05577_  (.A1(\soc/cpu/_01362_ ),
    .A2(\soc/cpu/_01370_ ),
    .B1(\soc/cpu/_01363_ ),
    .Y(\soc/cpu/_01371_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05578_  (.A1(\soc/cpu/_01116_ ),
    .A2(\soc/cpu/_01362_ ),
    .B1(\soc/cpu/_01371_ ),
    .B2(\soc/cpu/_01242_ ),
    .Y(\soc/cpu/_01372_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05579_  (.A(\soc/cpu/_01260_ ),
    .B(\soc/cpu/_01174_ ),
    .Y(\soc/cpu/_01373_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05580_  (.A1(\soc/cpu/_01181_ ),
    .A2(\soc/cpu/_01372_ ),
    .B1(\soc/cpu/_01373_ ),
    .Y(\soc/cpu/_01374_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05581_  (.A(\soc/cpu/_01160_ ),
    .B(\soc/cpu/_01374_ ),
    .Y(\soc/cpu/_01375_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05582_  (.A1(\soc/cpu/_01361_ ),
    .A2(\soc/cpu/_01370_ ),
    .B1(\soc/cpu/_01375_ ),
    .Y(\soc/cpu/_00047_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05583_  (.A1(\soc/cpu/_01050_ ),
    .A2(\soc/cpu/_01092_ ),
    .B1(\soc/cpu/_01090_ ),
    .B2(\soc/cpu/_01048_ ),
    .Y(\soc/cpu/_01376_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05584_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01376_ ),
    .B1(\soc/cpu/_01091_ ),
    .Y(\soc/cpu/_01377_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05585_  (.A(\soc/cpu/_01171_ ),
    .B(\soc/cpu/_01228_ ),
    .Y(\soc/cpu/_01378_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05586_  (.A(\soc/cpu/_01378_ ),
    .B(\soc/cpu/_01377_ ),
    .Y(\soc/cpu/_01379_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05587_  (.A(\soc/cpu/_01102_ ),
    .B(\soc/cpu/_01362_ ),
    .Y(\soc/cpu/_01380_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05588_  (.A(\soc/cpu/_01379_ ),
    .B(\soc/cpu/_01380_ ),
    .Y(\soc/cpu/_01381_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05589_  (.A1(\soc/cpu/_01363_ ),
    .A2(\soc/cpu/_01381_ ),
    .B1(\soc/cpu/_01181_ ),
    .Y(\soc/cpu/_01382_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_05590_  (.A1(\soc/cpu/_01166_ ),
    .A2(\soc/cpu/_01183_ ),
    .B1(\soc/cpu/_01358_ ),
    .B2(\soc/cpu/_01057_ ),
    .Y(\soc/cpu/_01383_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_05591_  (.A1(\soc/cpu/_01095_ ),
    .A2(\soc/cpu/_01235_ ),
    .A3(\soc/cpu/_01193_ ),
    .B1(\soc/cpu/_01383_ ),
    .B2(\soc/cpu/_01102_ ),
    .Y(\soc/cpu/_01384_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05592_  (.A1(\soc/cpu/_01367_ ),
    .A2(\soc/cpu/_01382_ ),
    .B1(\soc/cpu/_01384_ ),
    .Y(\soc/cpu/_01385_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05593_  (.A1(\soc/cpu/_01361_ ),
    .A2(\soc/cpu/_01377_ ),
    .B1(\soc/cpu/_01385_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00048_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_05594_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01143_ ),
    .B1(\soc/cpu/_01142_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01386_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05595_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01386_ ),
    .B1(\soc/cpu/_01141_ ),
    .Y(\soc/cpu/_01387_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05596_  (.A1(\soc/cpu/_01362_ ),
    .A2(\soc/cpu/_01387_ ),
    .B1(\soc/cpu/_01363_ ),
    .Y(\soc/cpu/_01388_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05597_  (.A1(\soc/cpu/_01210_ ),
    .A2(\soc/cpu/_01362_ ),
    .B1(\soc/cpu/_01388_ ),
    .Y(\soc/cpu/_01389_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05598_  (.A1(\soc/cpu/_01181_ ),
    .A2(\soc/cpu/_01389_ ),
    .B1(\soc/cpu/_01373_ ),
    .Y(\soc/cpu/_01390_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05599_  (.A(\soc/cpu/_01064_ ),
    .B(\soc/cpu/_01183_ ),
    .Y(\soc/cpu/_01391_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05600_  (.A1(\soc/cpu/_01235_ ),
    .A2(\soc/cpu/_01387_ ),
    .B1(\soc/cpu/_01193_ ),
    .Y(\soc/cpu/_01392_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/_05601_  (.A1(\soc/cpu/_01210_ ),
    .A2(\soc/cpu/_01211_ ),
    .B1(\soc/cpu/_01391_ ),
    .B2(\soc/cpu/_01228_ ),
    .C1(\soc/cpu/_01392_ ),
    .Y(\soc/cpu/_01393_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05602_  (.A1(\soc/cpu/_01088_ ),
    .A2(\soc/cpu/_01383_ ),
    .B1(\soc/cpu/_01393_ ),
    .Y(\soc/cpu/_01394_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05603_  (.A1(\soc/cpu/_01390_ ),
    .A2(\soc/cpu/_01394_ ),
    .B1(\soc/cpu/_01160_ ),
    .Y(\soc/cpu/_01395_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05604_  (.A1(\soc/cpu/_01360_ ),
    .A2(\soc/cpu/_01387_ ),
    .B1(\soc/cpu/_01395_ ),
    .Y(\soc/cpu/_00049_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_05605_  (.A1(\soc/cpu/_01048_ ),
    .A2(\soc/cpu/_01132_ ),
    .B1(\soc/cpu/_01135_ ),
    .B2(\soc/cpu/_01050_ ),
    .Y(\soc/cpu/_01396_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05606_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01396_ ),
    .B1(\soc/cpu/_01134_ ),
    .Y(\soc/cpu/_01397_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05607_  (.A(\soc/cpu/_01363_ ),
    .B(\soc/cpu/_01362_ ),
    .Y(\soc/cpu/_01398_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05608_  (.A1(\soc/cpu/_01226_ ),
    .A2(\soc/cpu/_01398_ ),
    .B1(\soc/cpu/_01289_ ),
    .Y(\soc/cpu/_01399_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05609_  (.A(\soc/cpu/_01363_ ),
    .B(\soc/cpu/_01378_ ),
    .C(\soc/cpu/_01397_ ),
    .Y(\soc/cpu/_01400_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05610_  (.A1(\soc/cpu/_01289_ ),
    .A2(\soc/cpu/_01183_ ),
    .B1(\soc/cpu/_01400_ ),
    .Y(\soc/cpu/_01401_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05611_  (.A1(\soc/cpu/_01181_ ),
    .A2(\soc/cpu/_01399_ ),
    .A3(\soc/cpu/_01401_ ),
    .B1(\soc/cpu/_01373_ ),
    .Y(\soc/cpu/_01402_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05612_  (.A(\soc/cpu/_01183_ ),
    .B(\soc/cpu/_01193_ ),
    .C(\soc/cpu/_01397_ ),
    .Y(\soc/cpu/_01403_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05613_  (.A(\soc/cpu/_01183_ ),
    .B(\soc/cpu/_01198_ ),
    .Y(\soc/cpu/_01404_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_05614_  (.A1(\soc/cpu/_01189_ ),
    .A2(\soc/cpu/_01095_ ),
    .A3(\soc/cpu/_01391_ ),
    .B1(\soc/cpu/_01404_ ),
    .B2(\soc/cpu/_01171_ ),
    .Y(\soc/cpu/_01405_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05615_  (.A(\soc/cpu/_01402_ ),
    .B(\soc/cpu/_01403_ ),
    .C(\soc/cpu/_01405_ ),
    .Y(\soc/cpu/_01406_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05616_  (.A1(\soc/cpu/_01360_ ),
    .A2(\soc/cpu/_01397_ ),
    .B1(\soc/cpu/_01406_ ),
    .B2(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_00050_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05617_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_01146_ ),
    .Y(\soc/cpu/_01407_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05618_  (.A1(\soc/cpu/mem_rdata_q[7] ),
    .A2(\soc/cpu/_00718_ ),
    .B1(\soc/cpu/_01407_ ),
    .Y(\soc/cpu/_01408_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05619_  (.A1(\soc/cpu/_01215_ ),
    .A2(\soc/cpu/_01286_ ),
    .B1(\soc/cpu/_01283_ ),
    .B2(\soc/cpu/_01408_ ),
    .Y(\soc/cpu/_00058_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_05620_  (.A_N(\soc/cpu/_00936_ ),
    .B(\soc/cpu/cpu_state[4] ),
    .Y(\soc/cpu/_01409_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05622_  (.A(\soc/cpu/cpuregs_raddr2[2] ),
    .Y(\soc/cpu/_01411_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05623_  (.A(\soc/cpu/cpuregs_raddr2[1] ),
    .B(\soc/cpu/cpuregs_raddr2[0] ),
    .Y(\soc/cpu/_01412_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_05624_  (.A(\soc/cpu/cpuregs_raddr2[3] ),
    .B(\soc/cpu/cpuregs_raddr2[2] ),
    .C(\soc/cpu/cpuregs_raddr2[4] ),
    .Y(\soc/cpu/_01413_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_05625_  (.A(\soc/cpu/_01412_ ),
    .B(\soc/cpu/_01413_ ),
    .Y(\soc/cpu/_01414_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05626_  (.A1(\soc/cpu/cpuregs_rdata2[2] ),
    .A2(\soc/cpu/_01414_ ),
    .B1(\soc/cpu/is_slli_srli_srai ),
    .Y(\soc/cpu/_01415_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/_05628_  (.A1(\soc/cpu/is_slli_srli_srai ),
    .A2(\soc/cpu/_01411_ ),
    .B1(\soc/cpu/_01415_ ),
    .C1(\soc/cpu/cpu_state[4] ),
    .X(\soc/cpu/_01417_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_05629_  (.A1(\soc/cpu/reg_sh[2] ),
    .A2(\soc/cpu/_01409_ ),
    .B1(\soc/cpu/_01417_ ),
    .C1(\soc/cpu/_00938_ ),
    .Y(\soc/cpu/_00061_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05631_  (.A1(\soc/cpu/cpuregs_rdata2[3] ),
    .A2(\soc/cpu/_01414_ ),
    .B1(\soc/cpu/is_slli_srli_srai ),
    .Y(\soc/cpu/_01419_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_05632_  (.A(\soc/cpu/is_slli_srli_srai ),
    .SLEEP(net963),
    .X(\soc/cpu/_01420_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_8 \soc/cpu/_05633_  (.A(\soc/cpu/cpu_state[4] ),
    .SLEEP(\soc/cpu/_00936_ ),
    .X(\soc/cpu/_01421_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05635_  (.A(\soc/cpu/reg_sh[2] ),
    .B(\soc/cpu/reg_sh[3] ),
    .Y(\soc/cpu/_01423_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05636_  (.A(\soc/cpu/_01421_ ),
    .B(\soc/cpu/_01423_ ),
    .Y(\soc/cpu/_01424_ ));
 sky130_fd_sc_hd__o311ai_1 \soc/cpu/_05637_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/_01419_ ),
    .A3(\soc/cpu/_01420_ ),
    .B1(\soc/cpu/_01424_ ),
    .C1(\soc/cpu/_00938_ ),
    .Y(\soc/cpu/_00062_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05638_  (.A1(\soc/cpu/reg_sh[2] ),
    .A2(\soc/cpu/reg_sh[3] ),
    .B1(\soc/cpu/reg_sh[4] ),
    .Y(\soc/cpu/_01425_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05639_  (.A(\soc/cpu/cpuregs_rdata2[4] ),
    .B(\soc/cpu/_01414_ ),
    .Y(\soc/cpu/_01426_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05640_  (.A(\soc/cpu/is_slli_srli_srai ),
    .B(\soc/cpu/_01426_ ),
    .Y(\soc/cpu/_01427_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_05641_  (.A1(\soc/cpu/is_slli_srli_srai ),
    .A2(net962),
    .B1(\soc/cpu/_01427_ ),
    .C1(\soc/cpu/cpu_state[4] ),
    .Y(\soc/cpu/_01428_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05642_  (.A1(\soc/cpu/_00979_ ),
    .A2(\soc/cpu/_01425_ ),
    .B1(\soc/cpu/_01428_ ),
    .Y(\soc/cpu/_00063_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_05643_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/cpu_state[5] ),
    .X(\soc/cpu/_01429_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05645_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(\soc/cpu/pcpi_rs2 [29]),
    .Y(\soc/cpu/_01431_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05646_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .B(\soc/cpu/pcpi_rs2 [28]),
    .Y(\soc/cpu/_01432_ ));
 sky130_fd_sc_hd__xor2_2 \soc/cpu/_05647_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .B(\soc/cpu/pcpi_rs2 [25]),
    .X(\soc/cpu/_01433_ ));
 sky130_fd_sc_hd__xnor2_4 \soc/cpu/_05649_  (.A(\soc/cpu/pcpi_rs1 [31]),
    .B(\soc/cpu/pcpi_rs2 [31]),
    .Y(\soc/cpu/_01435_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05651_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(\soc/cpu/pcpi_rs2 [30]),
    .Y(\soc/cpu/_01437_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05652_  (.A(\soc/cpu/_01435_ ),
    .B(\soc/cpu/_01437_ ),
    .Y(\soc/cpu/_01438_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05653_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(\soc/cpu/pcpi_rs2 [24]),
    .X(\soc/cpu/_01439_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05655_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(\soc/cpu/pcpi_rs2 [26]),
    .Y(\soc/cpu/_01441_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05656_  (.A(\soc/cpu/pcpi_rs1 [27]),
    .B(\soc/cpu/pcpi_rs2 [27]),
    .Y(\soc/cpu/_01442_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05657_  (.A(\soc/cpu/_01441_ ),
    .B(\soc/cpu/_01442_ ),
    .Y(\soc/cpu/_01443_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_05658_  (.A(\soc/cpu/_01433_ ),
    .B(\soc/cpu/_01438_ ),
    .C(\soc/cpu/_01439_ ),
    .D(\soc/cpu/_01443_ ),
    .Y(\soc/cpu/_01444_ ));
 sky130_fd_sc_hd__nand3_2 \soc/cpu/_05659_  (.A(\soc/cpu/_01431_ ),
    .B(\soc/cpu/_01432_ ),
    .C(\soc/cpu/_01444_ ),
    .Y(\soc/cpu/_01445_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05662_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(\soc/cpu/pcpi_rs2 [17]),
    .Y(\soc/cpu/_01448_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05665_  (.A(\soc/cpu/pcpi_rs1 [18]),
    .B(\soc/cpu/pcpi_rs2 [18]),
    .Y(\soc/cpu/_01451_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05667_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(\soc/cpu/pcpi_rs2 [16]),
    .Y(\soc/cpu/_01453_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_05668_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(\soc/cpu/pcpi_rs2 [19]),
    .Y(\soc/cpu/_01454_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_05669_  (.A(\soc/cpu/_01448_ ),
    .B(\soc/cpu/_01451_ ),
    .C(\soc/cpu/_01453_ ),
    .D(\soc/cpu/_01454_ ),
    .Y(\soc/cpu/_01455_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05670_  (.A(\soc/cpu/pcpi_rs1 [21]),
    .B(\soc/cpu/pcpi_rs2 [21]),
    .Y(\soc/cpu/_01456_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_05672_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(\soc/cpu/pcpi_rs2 [23]),
    .Y(\soc/cpu/_01458_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05674_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(net972),
    .Y(\soc/cpu/_01460_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05677_  (.A(\soc/cpu/pcpi_rs1 [20]),
    .B(\soc/cpu/pcpi_rs2 [20]),
    .Y(\soc/cpu/_01463_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_05678_  (.A(\soc/cpu/_01456_ ),
    .B(\soc/cpu/_01458_ ),
    .C(\soc/cpu/_01460_ ),
    .D(\soc/cpu/_01463_ ),
    .Y(\soc/cpu/_01464_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_05679_  (.A(\soc/cpu/_01445_ ),
    .B(\soc/cpu/_01455_ ),
    .C(\soc/cpu/_01464_ ),
    .Y(\soc/cpu/_01465_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05681_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/pcpi_rs2 [13]),
    .Y(\soc/cpu/_01467_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05684_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/pcpi_rs2 [12]),
    .Y(\soc/cpu/_01470_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05687_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(\soc/cpu/pcpi_rs2 [8]),
    .Y(\soc/cpu/_01473_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_05689_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(net781),
    .Y(\soc/cpu/_01475_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05690_  (.A(\soc/cpu/_01467_ ),
    .B(\soc/cpu/_01470_ ),
    .C(\soc/cpu/_01473_ ),
    .D(\soc/cpu/_01475_ ),
    .Y(\soc/cpu/_01476_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05692_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(\soc/cpu/pcpi_rs2 [15]),
    .Y(\soc/cpu/_01478_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05695_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(\soc/cpu/pcpi_rs2 [14]),
    .Y(\soc/cpu/_01481_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05696_  (.A(\soc/cpu/_01478_ ),
    .B(\soc/cpu/_01481_ ),
    .Y(\soc/cpu/_01482_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05698_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(\soc/cpu/pcpi_rs2 [11]),
    .Y(\soc/cpu/_01484_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05701_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(\soc/cpu/pcpi_rs2 [10]),
    .Y(\soc/cpu/_01487_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05702_  (.A(\soc/cpu/_01484_ ),
    .B(\soc/cpu/_01487_ ),
    .Y(\soc/cpu/_01488_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_05703_  (.A(\soc/cpu/_01476_ ),
    .B(\soc/cpu/_01482_ ),
    .C(\soc/cpu/_01488_ ),
    .Y(\soc/cpu/_01489_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05704_  (.A(\soc/cpu/pcpi_rs1 [0]),
    .Y(\soc/cpu/_01490_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05706_  (.A(\soc/cpu/_01490_ ),
    .B(\soc/cpu/mem_la_wdata [0]),
    .Y(\soc/cpu/_01492_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05707_  (.A(\soc/cpu/_01490_ ),
    .B(\soc/cpu/mem_la_wdata [0]),
    .Y(\soc/cpu/_01493_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_05708_  (.A(\soc/cpu/_01492_ ),
    .B_N(\soc/cpu/_01493_ ),
    .Y(\soc/cpu/_01494_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05710_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(\soc/cpu/mem_la_wdata [5]),
    .Y(\soc/cpu/_01496_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05712_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/mem_la_wdata [4]),
    .Y(\soc/cpu/_01498_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05714_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(net969),
    .Y(\soc/cpu/_01500_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_05715_  (.A(\soc/cpu/_01494_ ),
    .B(\soc/cpu/_01496_ ),
    .C(\soc/cpu/_01498_ ),
    .D(\soc/cpu/_01500_ ),
    .Y(\soc/cpu/_01501_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05717_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(\soc/cpu/mem_la_wdata [3]),
    .X(\soc/cpu/_01503_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05719_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/mem_la_wdata [2]),
    .Y(\soc/cpu/_01505_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_05720_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/mem_la_wdata [2]),
    .X(\soc/cpu/_01506_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05721_  (.A(\soc/cpu/_01505_ ),
    .B(\soc/cpu/_01506_ ),
    .Y(\soc/cpu/_01507_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05722_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(\soc/cpu/mem_la_wdata [7]),
    .Y(\soc/cpu/_01508_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05724_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(net776),
    .Y(\soc/cpu/_01510_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05725_  (.A(\soc/cpu/_01508_ ),
    .B(\soc/cpu/_01510_ ),
    .Y(\soc/cpu/_01511_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05726_  (.A(\soc/cpu/_01501_ ),
    .B(\soc/cpu/_01503_ ),
    .C(\soc/cpu/_01507_ ),
    .D(\soc/cpu/_01511_ ),
    .Y(\soc/cpu/_01512_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_05727_  (.A(\soc/cpu/_01465_ ),
    .B(\soc/cpu/_01489_ ),
    .C(\soc/cpu/_01512_ ),
    .Y(\soc/cpu/_01513_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_05728_  (.A(\soc/cpu/instr_bgeu ),
    .B(\soc/cpu/instr_bge ),
    .C(\soc/cpu/instr_bne ),
    .D(\soc/cpu/is_sltiu_bltu_sltu ),
    .X(\soc/cpu/_01514_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05729_  (.A(\soc/cpu/is_slti_blt_slt ),
    .B(\soc/cpu/_01514_ ),
    .Y(\soc/cpu/_01515_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05730_  (.A(net773),
    .Y(\soc/cpu/_01516_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05731_  (.A(\soc/cpu/mem_la_wdata [5]),
    .Y(\soc/cpu/_01517_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05732_  (.A(\soc/cpu/mem_la_wdata [4]),
    .Y(\soc/cpu/_01518_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05733_  (.A(\soc/cpu/mem_la_wdata [3]),
    .Y(\soc/cpu/_01519_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05734_  (.A(net855),
    .Y(\soc/cpu/_01520_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05735_  (.A(net848),
    .Y(\soc/cpu/_01521_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05736_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/_01521_ ),
    .C(\soc/cpu/_01492_ ),
    .X(\soc/cpu/_01522_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05737_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/_01520_ ),
    .C(\soc/cpu/_01522_ ),
    .X(\soc/cpu/_01523_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05738_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(\soc/cpu/_01519_ ),
    .C(\soc/cpu/_01523_ ),
    .X(\soc/cpu/_01524_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05739_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/_01518_ ),
    .C(\soc/cpu/_01524_ ),
    .X(\soc/cpu/_01525_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05740_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(\soc/cpu/_01517_ ),
    .C(\soc/cpu/_01525_ ),
    .X(\soc/cpu/_01526_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_05742_  (.A_N(\soc/cpu/pcpi_rs1 [6]),
    .B(\soc/cpu/mem_la_wdata [6]),
    .C(\soc/cpu/_01508_ ),
    .Y(\soc/cpu/_01528_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/_05743_  (.A1(\soc/cpu/pcpi_rs1 [7]),
    .A2(\soc/cpu/_01516_ ),
    .B1(\soc/cpu/_01511_ ),
    .B2(\soc/cpu/_01526_ ),
    .C1(\soc/cpu/_01528_ ),
    .Y(\soc/cpu/_01529_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05744_  (.A(\soc/cpu/pcpi_rs2 [15]),
    .Y(\soc/cpu/_01530_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05745_  (.A(\soc/cpu/pcpi_rs2 [14]),
    .B(\soc/cpu/_01478_ ),
    .Y(\soc/cpu/_01531_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05746_  (.A1(\soc/cpu/pcpi_rs1 [15]),
    .A2(\soc/cpu/_01530_ ),
    .B1(\soc/cpu/pcpi_rs1 [14]),
    .B2(\soc/cpu/_01531_ ),
    .Y(\soc/cpu/_01532_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05747_  (.A(\soc/cpu/pcpi_rs2 [13]),
    .Y(\soc/cpu/_01533_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05748_  (.A(\soc/cpu/pcpi_rs2 [12]),
    .Y(\soc/cpu/_01534_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05749_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .Y(\soc/cpu/_01535_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05751_  (.A(net777),
    .Y(\soc/cpu/_01537_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05752_  (.A(net781),
    .Y(\soc/cpu/_01538_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_05753_  (.A_N(\soc/cpu/pcpi_rs1 [8]),
    .B(\soc/cpu/pcpi_rs2 [8]),
    .C(\soc/cpu/_01475_ ),
    .Y(\soc/cpu/_01539_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05754_  (.A1(\soc/cpu/pcpi_rs1 [9]),
    .A2(\soc/cpu/_01538_ ),
    .B1(\soc/cpu/_01539_ ),
    .X(\soc/cpu/_01540_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_05755_  (.A1(\soc/cpu/pcpi_rs1 [11]),
    .A2(\soc/cpu/_01537_ ),
    .B1(\soc/cpu/_01488_ ),
    .B2(\soc/cpu/_01540_ ),
    .Y(\soc/cpu/_01541_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05756_  (.A1(\soc/cpu/_01535_ ),
    .A2(\soc/cpu/pcpi_rs2 [10]),
    .A3(\soc/cpu/_01484_ ),
    .B1(\soc/cpu/_01541_ ),
    .Y(\soc/cpu/_01542_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05757_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/_01534_ ),
    .C(\soc/cpu/_01542_ ),
    .X(\soc/cpu/_01543_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05758_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/_01533_ ),
    .C(\soc/cpu/_01543_ ),
    .X(\soc/cpu/_01544_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05759_  (.A(\soc/cpu/_01482_ ),
    .B(\soc/cpu/_01544_ ),
    .Y(\soc/cpu/_01545_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/_05760_  (.A1(\soc/cpu/_01489_ ),
    .A2(\soc/cpu/_01529_ ),
    .B1(\soc/cpu/_01532_ ),
    .C1(\soc/cpu/_01545_ ),
    .X(\soc/cpu/_01546_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05761_  (.A_N(\soc/cpu/pcpi_rs1 [23]),
    .B(\soc/cpu/pcpi_rs2 [23]),
    .Y(\soc/cpu/_01547_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_05763_  (.A_N(\soc/cpu/pcpi_rs1 [22]),
    .B(\soc/cpu/pcpi_rs2 [22]),
    .C(\soc/cpu/_01458_ ),
    .Y(\soc/cpu/_01549_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05765_  (.A(\soc/cpu/pcpi_rs2 [21]),
    .Y(\soc/cpu/_01551_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05766_  (.A(\soc/cpu/pcpi_rs1 [20]),
    .Y(\soc/cpu/_01552_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05768_  (.A(\soc/cpu/pcpi_rs2 [19]),
    .Y(\soc/cpu/_01554_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05769_  (.A(\soc/cpu/pcpi_rs1 [18]),
    .Y(\soc/cpu/_01555_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_05770_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .Y(\soc/cpu/_01556_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_05771_  (.A(\soc/cpu/pcpi_rs2 [16]),
    .SLEEP(\soc/cpu/pcpi_rs1 [16]),
    .X(\soc/cpu/_01557_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05772_  (.A(\soc/cpu/_01556_ ),
    .B(\soc/cpu/pcpi_rs2 [17]),
    .C(\soc/cpu/_01557_ ),
    .X(\soc/cpu/_01558_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05773_  (.A(\soc/cpu/_01555_ ),
    .B(\soc/cpu/pcpi_rs2 [18]),
    .C(\soc/cpu/_01558_ ),
    .X(\soc/cpu/_01559_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05774_  (.A(\soc/cpu/_01454_ ),
    .B(\soc/cpu/_01559_ ),
    .Y(\soc/cpu/_01560_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05775_  (.A1(\soc/cpu/pcpi_rs1 [19]),
    .A2(\soc/cpu/_01554_ ),
    .B1(\soc/cpu/_01560_ ),
    .Y(\soc/cpu/_01561_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05776_  (.A(\soc/cpu/_01552_ ),
    .B(\soc/cpu/pcpi_rs2 [20]),
    .C(\soc/cpu/_01561_ ),
    .X(\soc/cpu/_01562_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05777_  (.A(\soc/cpu/_01456_ ),
    .B(\soc/cpu/_01562_ ),
    .Y(\soc/cpu/_01563_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05778_  (.A1(\soc/cpu/pcpi_rs1 [21]),
    .A2(\soc/cpu/_01551_ ),
    .B1(\soc/cpu/_01563_ ),
    .Y(\soc/cpu/_01564_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05779_  (.A(\soc/cpu/_01458_ ),
    .B(\soc/cpu/_01460_ ),
    .C(\soc/cpu/_01564_ ),
    .Y(\soc/cpu/_01565_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_05780_  (.A1(\soc/cpu/_01547_ ),
    .A2(\soc/cpu/_01549_ ),
    .A3(\soc/cpu/_01565_ ),
    .B1(\soc/cpu/_01445_ ),
    .Y(\soc/cpu/_01566_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05781_  (.A(\soc/cpu/pcpi_rs2 [29]),
    .Y(\soc/cpu/_01567_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05782_  (.A(\soc/cpu/pcpi_rs2 [28]),
    .Y(\soc/cpu/_01568_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05783_  (.A(\soc/cpu/pcpi_rs2 [27]),
    .Y(\soc/cpu/_01569_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05784_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .Y(\soc/cpu/_01570_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/cpu/_05785_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(\soc/cpu/_01433_ ),
    .C_N(\soc/cpu/pcpi_rs2 [24]),
    .Y(\soc/cpu/_01571_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05786_  (.A1(\soc/cpu/_01570_ ),
    .A2(\soc/cpu/pcpi_rs2 [25]),
    .B1(\soc/cpu/_01571_ ),
    .Y(\soc/cpu/_01572_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_05787_  (.A_N(\soc/cpu/pcpi_rs1 [26]),
    .B(\soc/cpu/pcpi_rs2 [26]),
    .C(\soc/cpu/_01442_ ),
    .Y(\soc/cpu/_01573_ ));
 sky130_fd_sc_hd__o221a_1 \soc/cpu/_05788_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(\soc/cpu/_01569_ ),
    .B1(\soc/cpu/_01443_ ),
    .B2(\soc/cpu/_01572_ ),
    .C1(\soc/cpu/_01573_ ),
    .X(\soc/cpu/_01574_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_05789_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .B(\soc/cpu/_01568_ ),
    .C(\soc/cpu/_01574_ ),
    .X(\soc/cpu/_01575_ ));
 sky130_fd_sc_hd__maj3_2 \soc/cpu/_05790_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(\soc/cpu/_01567_ ),
    .C(\soc/cpu/_01575_ ),
    .X(\soc/cpu/_01576_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05791_  (.A(\soc/cpu/pcpi_rs2 [30]),
    .B(\soc/cpu/_01435_ ),
    .Y(\soc/cpu/_01577_ ));
 sky130_fd_sc_hd__nand2b_2 \soc/cpu/_05792_  (.A_N(\soc/cpu/pcpi_rs1 [31]),
    .B(\soc/cpu/pcpi_rs2 [31]),
    .Y(\soc/cpu/_01578_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/_05793_  (.A1(\soc/cpu/_01438_ ),
    .A2(\soc/cpu/_01576_ ),
    .B1(\soc/cpu/_01577_ ),
    .B2(\soc/cpu/pcpi_rs1 [30]),
    .C1(\soc/cpu/_01578_ ),
    .Y(\soc/cpu/_01579_ ));
 sky130_fd_sc_hd__a211o_4 \soc/cpu/_05794_  (.A1(\soc/cpu/_01465_ ),
    .A2(\soc/cpu/_01546_ ),
    .B1(\soc/cpu/_01566_ ),
    .C1(\soc/cpu/_01579_ ),
    .X(\soc/cpu/_01580_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_05795_  (.A1(\soc/cpu/is_sltiu_bltu_sltu ),
    .A2(\soc/cpu/_01513_ ),
    .A3(\soc/cpu/_01580_ ),
    .B1(\soc/cpu/_01515_ ),
    .Y(\soc/cpu/_01581_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05796_  (.A(\soc/cpu/_01513_ ),
    .B(\soc/cpu/_01580_ ),
    .Y(\soc/cpu/_01582_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05797_  (.A_N(\soc/cpu/_01580_ ),
    .B(\soc/cpu/_01435_ ),
    .Y(\soc/cpu/_01583_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_05798_  (.A(\soc/cpu/_01513_ ),
    .B(\soc/cpu/_01578_ ),
    .C(\soc/cpu/_01583_ ),
    .Y(\soc/cpu/_01584_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_05799_  (.A0(\soc/cpu/is_slti_blt_slt ),
    .A1(\soc/cpu/instr_bge ),
    .S(\soc/cpu/_01584_ ),
    .X(\soc/cpu/_01585_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_05800_  (.A1(\soc/cpu/instr_bne ),
    .A2(\soc/cpu/_01513_ ),
    .B1(\soc/cpu/_01582_ ),
    .B2(\soc/cpu/instr_bgeu ),
    .C1(\soc/cpu/_01585_ ),
    .Y(\soc/cpu/_01586_ ));
 sky130_fd_sc_hd__a22o_4 \soc/cpu/_05801_  (.A1(\soc/cpu/_01513_ ),
    .A2(\soc/cpu/_01515_ ),
    .B1(\soc/cpu/_01581_ ),
    .B2(\soc/cpu/_01586_ ),
    .X(\soc/cpu/_01587_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_16 \soc/cpu/_05802_  (.A(\soc/cpu/mem_do_rinst ),
    .SLEEP(\soc/cpu/_00833_ ),
    .X(\soc/cpu/_01588_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05804_  (.A(\soc/cpu/mem_do_prefetch ),
    .B(\soc/cpu/_00833_ ),
    .C(\soc/cpu/_00838_ ),
    .Y(\soc/cpu/_00174_ ));
 sky130_fd_sc_hd__o32a_1 \soc/cpu/_05805_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_00917_ ),
    .A3(\soc/cpu/_01587_ ),
    .B1(\soc/cpu/_01588_ ),
    .B2(\soc/cpu/_00174_ ),
    .X(\soc/cpu/_00000_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05806_  (.A1(\soc/cpu/_01050_ ),
    .A2(\soc/cpu/_01075_ ),
    .B1(\soc/cpu/_01073_ ),
    .B2(\soc/cpu/_01048_ ),
    .Y(\soc/cpu/_01590_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_05807_  (.A1(\soc/cpu/_00718_ ),
    .A2(\soc/cpu/_01590_ ),
    .B1(\soc/cpu/_01074_ ),
    .Y(\soc/cpu/_01591_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05808_  (.A(\soc/cpu/_01165_ ),
    .B(\soc/cpu/_01264_ ),
    .Y(\soc/cpu/_01592_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05809_  (.A1(\soc/cpu/_01178_ ),
    .A2(\soc/cpu/_01592_ ),
    .B1(\soc/cpu/_01166_ ),
    .Y(\soc/cpu/_01593_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05810_  (.A(\soc/cpu/_01331_ ),
    .B(\soc/cpu/_01240_ ),
    .C(\soc/cpu/_01593_ ),
    .Y(\soc/cpu/_01594_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05811_  (.A1(\soc/cpu/_01266_ ),
    .A2(\soc/cpu/_01591_ ),
    .B1(\soc/cpu/_01201_ ),
    .Y(\soc/cpu/_01595_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05812_  (.A(\soc/cpu/_01594_ ),
    .B(\soc/cpu/_01595_ ),
    .Y(\soc/cpu/_01596_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05813_  (.A1(\soc/cpu/_01303_ ),
    .A2(\soc/cpu/_01591_ ),
    .B1(\soc/cpu/_01596_ ),
    .Y(\soc/cpu/_00057_ ));
 sky130_fd_sc_hd__a21o_2 \soc/cpu/_05814_  (.A1(\soc/cpu/latched_store ),
    .A2(\soc/cpu/latched_branch ),
    .B1(\soc/cpu/reg_next_pc[2] ),
    .X(\soc/cpu/_01597_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05815_  (.A1(\soc/cpu/reg_out[2] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01597_ ),
    .Y(\soc/cpu/_01598_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05816_  (.A(\soc/cpu/_00741_ ),
    .B(\soc/cpu/_01598_ ),
    .Y(\soc/cpu/_01599_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05818_  (.A(\soc/cpu/_00741_ ),
    .B(\soc/cpu/_01598_ ),
    .Y(\soc/cpu/_01601_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05819_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_01601_ ),
    .Y(\soc/cpu/_01602_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05821_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01604_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05822_  (.A1(\soc/cpu/_01599_ ),
    .A2(\soc/cpu/_01602_ ),
    .B1(\soc/cpu/_01604_ ),
    .Y(\soc/cpu/mem_la_addr [2]));
 sky130_fd_sc_hd__a21o_2 \soc/cpu/_05824_  (.A1(\soc/cpu/latched_store ),
    .A2(\soc/cpu/latched_branch ),
    .B1(\soc/cpu/reg_next_pc[3] ),
    .X(\soc/cpu/_01606_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05825_  (.A1(\soc/cpu/reg_out[3] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01606_ ),
    .Y(\soc/cpu/_01607_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05826_  (.A(\soc/cpu/_01599_ ),
    .B(\soc/cpu/_01607_ ),
    .X(\soc/cpu/_01608_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05827_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01609_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05828_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_01608_ ),
    .B1(\soc/cpu/_01609_ ),
    .Y(\soc/cpu/mem_la_addr [3]));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_05829_  (.A(\soc/cpu/_00741_ ),
    .B(\soc/cpu/_01598_ ),
    .C(\soc/cpu/_01607_ ),
    .X(\soc/cpu/_01610_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05830_  (.A0(\soc/cpu/reg_out[4] ),
    .A1(\soc/cpu/reg_next_pc[4] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01611_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05831_  (.A(\soc/cpu/_01610_ ),
    .B(\soc/cpu/_01611_ ),
    .Y(\soc/cpu/_01612_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_05833_  (.A1(\soc/cpu/_01610_ ),
    .A2(\soc/cpu/_01611_ ),
    .B1(\soc/cpu/_01159_ ),
    .X(\soc/cpu/_01614_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05835_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01616_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05836_  (.A1(\soc/cpu/_01612_ ),
    .A2(\soc/cpu/_01614_ ),
    .B1(\soc/cpu/_01616_ ),
    .Y(\soc/cpu/mem_la_addr [4]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05838_  (.A0(\soc/cpu/reg_out[5] ),
    .A1(\soc/cpu/reg_next_pc[5] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01618_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05839_  (.A(\soc/cpu/_01612_ ),
    .B(\soc/cpu/_01618_ ),
    .X(\soc/cpu/_01619_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05840_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01620_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05841_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_01619_ ),
    .B1(\soc/cpu/_01620_ ),
    .Y(\soc/cpu/mem_la_addr [5]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05843_  (.A0(\soc/cpu/reg_out[6] ),
    .A1(\soc/cpu/reg_next_pc[6] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01622_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05844_  (.A(\soc/cpu/_01610_ ),
    .B(\soc/cpu/_01611_ ),
    .C(\soc/cpu/_01618_ ),
    .D(\soc/cpu/_01622_ ),
    .Y(\soc/cpu/_01623_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_05845_  (.A1(\soc/cpu/_01610_ ),
    .A2(\soc/cpu/_01611_ ),
    .A3(\soc/cpu/_01618_ ),
    .B1(\soc/cpu/_01622_ ),
    .Y(\soc/cpu/_01624_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05846_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_01624_ ),
    .Y(\soc/cpu/_01625_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05847_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01626_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05848_  (.A1(\soc/cpu/_01623_ ),
    .A2(\soc/cpu/_01625_ ),
    .B1(\soc/cpu/_01626_ ),
    .Y(\soc/cpu/mem_la_addr [6]));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_05850_  (.A(\soc/cpu/reg_next_pc[7] ),
    .B(net161),
    .Y(\soc/cpu/_01628_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05851_  (.A(\soc/cpu/reg_out[7] ),
    .B(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01629_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05852_  (.A(\soc/cpu/_01628_ ),
    .B(\soc/cpu/_01629_ ),
    .Y(\soc/cpu/_01630_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05853_  (.A(\soc/cpu/_01623_ ),
    .B(\soc/cpu/_01630_ ),
    .Y(\soc/cpu/_01631_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05855_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01633_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05856_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_01631_ ),
    .B1(\soc/cpu/_01633_ ),
    .Y(\soc/cpu/mem_la_addr [7]));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05857_  (.A0(\soc/cpu/reg_out[8] ),
    .A1(\soc/cpu/reg_next_pc[8] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01634_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05858_  (.A(\soc/cpu/_01634_ ),
    .Y(\soc/cpu/_01635_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05859_  (.A(\soc/cpu/_01623_ ),
    .B(\soc/cpu/_01630_ ),
    .C(\soc/cpu/_01635_ ),
    .Y(\soc/cpu/_01636_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05860_  (.A1(\soc/cpu/_01623_ ),
    .A2(\soc/cpu/_01630_ ),
    .B1(\soc/cpu/_01635_ ),
    .Y(\soc/cpu/_01637_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05861_  (.A(\soc/cpu/_01159_ ),
    .B(\soc/cpu/_01637_ ),
    .Y(\soc/cpu/_01638_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_05862_  (.A1(\soc/cpu/pcpi_rs1 [8]),
    .A2(\soc/cpu/_01159_ ),
    .B1(\soc/cpu/_01636_ ),
    .B2(\soc/cpu/_01638_ ),
    .X(\soc/cpu/mem_la_addr [8]));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05863_  (.A(\soc/cpu/reg_next_pc[9] ),
    .B(net161),
    .Y(\soc/cpu/_01639_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_05864_  (.A1(\soc/cpu/reg_out[9] ),
    .A2(\soc/cpu/_00709_ ),
    .B1_N(\soc/cpu/_01639_ ),
    .Y(\soc/cpu/_01640_ ));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_05865_  (.A(\soc/cpu/_01636_ ),
    .B(\soc/cpu/_01640_ ),
    .X(\soc/cpu/_01641_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05867_  (.A1(\soc/cpu/_01636_ ),
    .A2(\soc/cpu/_01640_ ),
    .B1(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01643_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_05868_  (.A1(\soc/cpu/pcpi_rs1 [9]),
    .A2(\soc/cpu/_01159_ ),
    .B1(\soc/cpu/_01641_ ),
    .B2(\soc/cpu/_01643_ ),
    .X(\soc/cpu/mem_la_addr [9]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05869_  (.A0(\soc/cpu/reg_out[10] ),
    .A1(\soc/cpu/reg_next_pc[10] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01644_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05870_  (.A(\soc/cpu/_01641_ ),
    .B(\soc/cpu/_01644_ ),
    .Y(\soc/cpu/_01645_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05871_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01646_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05872_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_01645_ ),
    .B1(\soc/cpu/_01646_ ),
    .Y(\soc/cpu/mem_la_addr [10]));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05873_  (.A(\soc/cpu/_01641_ ),
    .B(\soc/cpu/_01644_ ),
    .Y(\soc/cpu/_01647_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05874_  (.A0(\soc/cpu/reg_out[11] ),
    .A1(\soc/cpu/reg_next_pc[11] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01648_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05875_  (.A(\soc/cpu/_01647_ ),
    .B(\soc/cpu/_01648_ ),
    .X(\soc/cpu/_01649_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05877_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01651_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05878_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_01649_ ),
    .B1(\soc/cpu/_01651_ ),
    .Y(\soc/cpu/mem_la_addr [11]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05880_  (.A0(\soc/cpu/reg_out[12] ),
    .A1(\soc/cpu/reg_next_pc[12] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01653_ ));
 sky130_fd_sc_hd__nor4_4 \soc/cpu/_05881_  (.A(\soc/cpu/_01641_ ),
    .B(\soc/cpu/_01644_ ),
    .C(\soc/cpu/_01648_ ),
    .D(\soc/cpu/_01653_ ),
    .Y(\soc/cpu/_01654_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_05882_  (.A1(\soc/cpu/_01641_ ),
    .A2(\soc/cpu/_01644_ ),
    .A3(\soc/cpu/_01648_ ),
    .B1(\soc/cpu/_01653_ ),
    .Y(\soc/cpu/_01655_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05883_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_01655_ ),
    .Y(\soc/cpu/_01656_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05884_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01657_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05885_  (.A1(\soc/cpu/_01654_ ),
    .A2(\soc/cpu/_01656_ ),
    .B1(\soc/cpu/_01657_ ),
    .Y(\soc/cpu/mem_la_addr [12]));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_05887_  (.A(\soc/cpu/reg_next_pc[13] ),
    .B(net161),
    .X(\soc/cpu/_01659_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_05888_  (.A1(\soc/cpu/reg_out[13] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01659_ ),
    .X(\soc/cpu/_01660_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05889_  (.A(\soc/cpu/_01654_ ),
    .B(\soc/cpu/_01660_ ),
    .Y(\soc/cpu/_01661_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05890_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/_01159_ ),
    .Y(\soc/cpu/_01662_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05891_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_01661_ ),
    .B1(\soc/cpu/_01662_ ),
    .Y(\soc/cpu/mem_la_addr [13]));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05892_  (.A0(\soc/cpu/reg_out[14] ),
    .A1(\soc/cpu/reg_next_pc[14] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01663_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05893_  (.A(\soc/cpu/_01663_ ),
    .Y(\soc/cpu/_01664_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_05894_  (.A(\soc/cpu/_01654_ ),
    .B(\soc/cpu/_01660_ ),
    .C(\soc/cpu/_01664_ ),
    .Y(\soc/cpu/_01665_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05895_  (.A1(\soc/cpu/_01654_ ),
    .A2(\soc/cpu/_01660_ ),
    .B1(\soc/cpu/_01664_ ),
    .Y(\soc/cpu/_01666_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05896_  (.A(net158),
    .B(\soc/cpu/_01666_ ),
    .Y(\soc/cpu/_01667_ ));
 sky130_fd_sc_hd__a22o_2 \soc/cpu/_05897_  (.A1(\soc/cpu/pcpi_rs1 [14]),
    .A2(net158),
    .B1(\soc/cpu/_01665_ ),
    .B2(\soc/cpu/_01667_ ),
    .X(\soc/cpu/mem_la_addr [14]));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05898_  (.A0(\soc/cpu/reg_out[15] ),
    .A1(\soc/cpu/reg_next_pc[15] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01668_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_05899_  (.A(\soc/cpu/_01665_ ),
    .B(\soc/cpu/_01668_ ),
    .X(\soc/cpu/_01669_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05900_  (.A1(\soc/cpu/_01665_ ),
    .A2(\soc/cpu/_01668_ ),
    .B1(net158),
    .Y(\soc/cpu/_01670_ ));
 sky130_fd_sc_hd__a22o_2 \soc/cpu/_05901_  (.A1(\soc/cpu/pcpi_rs1 [15]),
    .A2(net158),
    .B1(\soc/cpu/_01669_ ),
    .B2(\soc/cpu/_01670_ ),
    .X(\soc/cpu/mem_la_addr [15]));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05902_  (.A0(\soc/cpu/reg_out[16] ),
    .A1(\soc/cpu/reg_next_pc[16] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01671_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_05903_  (.A(\soc/cpu/_01669_ ),
    .B(\soc/cpu/_01671_ ),
    .Y(\soc/cpu/_01672_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05904_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(net158),
    .Y(\soc/cpu/_01673_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05905_  (.A1(net158),
    .A2(\soc/cpu/_01672_ ),
    .B1(\soc/cpu/_01673_ ),
    .Y(\soc/cpu/mem_la_addr [16]));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_05906_  (.A0(\soc/cpu/reg_out[17] ),
    .A1(\soc/cpu/reg_next_pc[17] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01674_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05907_  (.A1(\soc/cpu/_01669_ ),
    .A2(\soc/cpu/_01671_ ),
    .B1(\soc/cpu/_01674_ ),
    .Y(\soc/cpu/_01675_ ));
 sky130_fd_sc_hd__or3_2 \soc/cpu/_05908_  (.A(\soc/cpu/_01669_ ),
    .B(\soc/cpu/_01671_ ),
    .C(\soc/cpu/_01674_ ),
    .X(\soc/cpu/_01676_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_05909_  (.A1(\soc/cpu/_01675_ ),
    .A2(\soc/cpu/_01676_ ),
    .B1(net158),
    .Y(\soc/cpu/_01677_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_05910_  (.A1(\soc/cpu/_01556_ ),
    .A2(net158),
    .B1(\soc/cpu/_01677_ ),
    .Y(\soc/cpu/mem_la_addr [17]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05912_  (.A0(\soc/cpu/reg_out[18] ),
    .A1(\soc/cpu/reg_next_pc[18] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01679_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05913_  (.A(\soc/cpu/_01676_ ),
    .B(\soc/cpu/_01679_ ),
    .Y(\soc/cpu/_01680_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_05914_  (.A1(\soc/cpu/_01676_ ),
    .A2(\soc/cpu/_01679_ ),
    .B1(net158),
    .X(\soc/cpu/_01681_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05915_  (.A1(\soc/cpu/_01555_ ),
    .A2(\soc/cpu/_00711_ ),
    .B1(\soc/cpu/_01680_ ),
    .B2(\soc/cpu/_01681_ ),
    .Y(\soc/cpu/mem_la_addr [18]));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_05917_  (.A(\soc/cpu/reg_next_pc[19] ),
    .B(\soc/cpu/_00707_ ),
    .X(\soc/cpu/_01683_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_05918_  (.A1(\soc/cpu/reg_out[19] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01683_ ),
    .Y(\soc/cpu/_01684_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05919_  (.A(\soc/cpu/_01680_ ),
    .B(\soc/cpu/_01684_ ),
    .X(\soc/cpu/_01685_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05920_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(net158),
    .Y(\soc/cpu/_01686_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05921_  (.A1(net158),
    .A2(\soc/cpu/_01685_ ),
    .B1(\soc/cpu/_01686_ ),
    .Y(\soc/cpu/mem_la_addr [19]));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05922_  (.A0(\soc/cpu/reg_out[20] ),
    .A1(\soc/cpu/reg_next_pc[20] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01687_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_05923_  (.A(\soc/cpu/_01676_ ),
    .B(\soc/cpu/_01679_ ),
    .C(\soc/cpu/_01684_ ),
    .D(\soc/cpu/_01687_ ),
    .Y(\soc/cpu/_01688_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05924_  (.A(\soc/cpu/_01676_ ),
    .B(\soc/cpu/_01679_ ),
    .C(\soc/cpu/_01684_ ),
    .Y(\soc/cpu/_01689_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_05925_  (.A_N(\soc/cpu/_01689_ ),
    .B(\soc/cpu/_01687_ ),
    .Y(\soc/cpu/_01690_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05926_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_01690_ ),
    .Y(\soc/cpu/_01691_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_05927_  (.A1(\soc/cpu/_01552_ ),
    .A2(\soc/cpu/_00711_ ),
    .B1(\soc/cpu/_01688_ ),
    .B2(\soc/cpu/_01691_ ),
    .Y(\soc/cpu/mem_la_addr [20]));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_05929_  (.A(\soc/cpu/reg_next_pc[21] ),
    .B(\soc/cpu/_00707_ ),
    .X(\soc/cpu/_01693_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05930_  (.A1(\soc/cpu/reg_out[21] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01693_ ),
    .Y(\soc/cpu/_01694_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05931_  (.A(\soc/cpu/_01688_ ),
    .B(\soc/cpu/_01694_ ),
    .X(\soc/cpu/_01695_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05932_  (.A(\soc/cpu/pcpi_rs1 [21]),
    .B(net158),
    .Y(\soc/cpu/_01696_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05933_  (.A1(net158),
    .A2(\soc/cpu/_01695_ ),
    .B1(\soc/cpu/_01696_ ),
    .Y(\soc/cpu/mem_la_addr [21]));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_05934_  (.A(\soc/cpu/_01688_ ),
    .SLEEP(\soc/cpu/_01694_ ),
    .X(\soc/cpu/_01697_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_05936_  (.A(\soc/cpu/reg_next_pc[22] ),
    .B(\soc/cpu/_00707_ ),
    .X(\soc/cpu/_01699_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_05937_  (.A1(\soc/cpu/reg_out[22] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01699_ ),
    .Y(\soc/cpu/_01700_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05938_  (.A(\soc/cpu/_01697_ ),
    .B(\soc/cpu/_01700_ ),
    .X(\soc/cpu/_01701_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05939_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(net158),
    .Y(\soc/cpu/_01702_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05940_  (.A1(net158),
    .A2(\soc/cpu/_01701_ ),
    .B1(\soc/cpu/_01702_ ),
    .Y(\soc/cpu/mem_la_addr [22]));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_05941_  (.A1(\soc/cpu/reg_out[22] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01697_ ),
    .C1(\soc/cpu/_01699_ ),
    .Y(\soc/cpu/_01703_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05942_  (.A0(\soc/cpu/reg_out[23] ),
    .A1(\soc/cpu/reg_next_pc[23] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01704_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05943_  (.A(\soc/cpu/_01703_ ),
    .B(\soc/cpu/_01704_ ),
    .Y(\soc/cpu/_01705_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_05944_  (.A1(\soc/cpu/_01703_ ),
    .A2(\soc/cpu/_01704_ ),
    .B1(net158),
    .X(\soc/cpu/_01706_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05946_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(net158),
    .Y(\soc/cpu/_01708_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05947_  (.A1(\soc/cpu/_01705_ ),
    .A2(\soc/cpu/_01706_ ),
    .B1(\soc/cpu/_01708_ ),
    .Y(\soc/cpu/mem_la_addr [23]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05948_  (.A0(\soc/cpu/reg_out[24] ),
    .A1(\soc/cpu/reg_next_pc[24] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01709_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05949_  (.A(\soc/cpu/_01705_ ),
    .B(\soc/cpu/_01709_ ),
    .X(\soc/cpu/_01710_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05951_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(net158),
    .Y(\soc/cpu/_01712_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05952_  (.A1(net158),
    .A2(\soc/cpu/_01710_ ),
    .B1(\soc/cpu/_01712_ ),
    .Y(\soc/cpu/mem_la_addr [24]));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05953_  (.A(\soc/cpu/_01703_ ),
    .B(\soc/cpu/_01704_ ),
    .C(\soc/cpu/_01709_ ),
    .Y(\soc/cpu/_01713_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05954_  (.A0(\soc/cpu/reg_out[25] ),
    .A1(\soc/cpu/reg_next_pc[25] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01714_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05955_  (.A(\soc/cpu/_01713_ ),
    .B(\soc/cpu/_01714_ ),
    .X(\soc/cpu/_01715_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05957_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .B(net158),
    .Y(\soc/cpu/_01717_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05958_  (.A1(net158),
    .A2(\soc/cpu/_01715_ ),
    .B1(\soc/cpu/_01717_ ),
    .Y(\soc/cpu/mem_la_addr [25]));
 sky130_fd_sc_hd__or4_2 \soc/cpu/_05959_  (.A(\soc/cpu/_01703_ ),
    .B(\soc/cpu/_01704_ ),
    .C(\soc/cpu/_01709_ ),
    .D(\soc/cpu/_01714_ ),
    .X(\soc/cpu/_01718_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05960_  (.A0(\soc/cpu/reg_out[26] ),
    .A1(\soc/cpu/reg_next_pc[26] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01719_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05961_  (.A(\soc/cpu/_01718_ ),
    .B(\soc/cpu/_01719_ ),
    .Y(\soc/cpu/_01720_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05962_  (.A(\soc/cpu/_01718_ ),
    .B(\soc/cpu/_01719_ ),
    .Y(\soc/cpu/_01721_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05963_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_01721_ ),
    .Y(\soc/cpu/_01722_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05965_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(net158),
    .Y(\soc/cpu/_01724_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05966_  (.A1(\soc/cpu/_01720_ ),
    .A2(\soc/cpu/_01722_ ),
    .B1(\soc/cpu/_01724_ ),
    .Y(\soc/cpu/mem_la_addr [26]));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05967_  (.A0(\soc/cpu/reg_out[27] ),
    .A1(\soc/cpu/reg_next_pc[27] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01725_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05968_  (.A(\soc/cpu/_01720_ ),
    .B(\soc/cpu/_01725_ ),
    .X(\soc/cpu/_01726_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05970_  (.A(\soc/cpu/pcpi_rs1 [27]),
    .B(net158),
    .Y(\soc/cpu/_01728_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05971_  (.A1(net158),
    .A2(\soc/cpu/_01726_ ),
    .B1(\soc/cpu/_01728_ ),
    .Y(\soc/cpu/mem_la_addr [27]));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05972_  (.A(\soc/cpu/_01718_ ),
    .B(\soc/cpu/_01719_ ),
    .C(\soc/cpu/_01725_ ),
    .Y(\soc/cpu/_01729_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_05974_  (.A(\soc/cpu/reg_next_pc[28] ),
    .B(\soc/cpu/_00707_ ),
    .X(\soc/cpu/_01731_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_05975_  (.A1(\soc/cpu/reg_out[28] ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_01731_ ),
    .Y(\soc/cpu/_01732_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05976_  (.A(\soc/cpu/_01729_ ),
    .B(\soc/cpu/_01732_ ),
    .X(\soc/cpu/_01733_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05978_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .B(net158),
    .Y(\soc/cpu/_01735_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05979_  (.A1(net158),
    .A2(\soc/cpu/_01733_ ),
    .B1(\soc/cpu/_01735_ ),
    .Y(\soc/cpu/mem_la_addr [28]));
 sky130_fd_sc_hd__or4_2 \soc/cpu/_05980_  (.A(\soc/cpu/_01718_ ),
    .B(\soc/cpu/_01719_ ),
    .C(\soc/cpu/_01725_ ),
    .D(\soc/cpu/_01732_ ),
    .X(\soc/cpu/_01736_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05981_  (.A0(\soc/cpu/reg_out[29] ),
    .A1(\soc/cpu/reg_next_pc[29] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01737_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05982_  (.A(\soc/cpu/_01736_ ),
    .B(\soc/cpu/_01737_ ),
    .Y(\soc/cpu/_01738_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05983_  (.A(\soc/cpu/_01736_ ),
    .B(\soc/cpu/_01737_ ),
    .Y(\soc/cpu/_01739_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05984_  (.A(\soc/cpu/_00711_ ),
    .B(\soc/cpu/_01739_ ),
    .Y(\soc/cpu/_01740_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_05986_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(net158),
    .Y(\soc/cpu/_01742_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05987_  (.A1(\soc/cpu/_01738_ ),
    .A2(\soc/cpu/_01740_ ),
    .B1(\soc/cpu/_01742_ ),
    .Y(\soc/cpu/mem_la_addr [29]));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_05988_  (.A0(\soc/cpu/reg_out[30] ),
    .A1(\soc/cpu/reg_next_pc[30] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01743_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05989_  (.A(\soc/cpu/_01738_ ),
    .B(\soc/cpu/_01743_ ),
    .X(\soc/cpu/_01744_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_05991_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(net158),
    .Y(\soc/cpu/_01746_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_05992_  (.A1(net158),
    .A2(\soc/cpu/_01744_ ),
    .B1(\soc/cpu/_01746_ ),
    .Y(\soc/cpu/mem_la_addr [30]));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_05993_  (.A(\soc/cpu/_01736_ ),
    .B(\soc/cpu/_01737_ ),
    .C(\soc/cpu/_01743_ ),
    .Y(\soc/cpu/_01747_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_05994_  (.A0(\soc/cpu/reg_out[31] ),
    .A1(\soc/cpu/reg_next_pc[31] ),
    .S(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_01748_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_05995_  (.A(\soc/cpu/_01747_ ),
    .B(\soc/cpu/_01748_ ),
    .X(\soc/cpu/_01749_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_05996_  (.A(\soc/cpu/pcpi_rs1 [31]),
    .B(\soc/cpu/_00711_ ),
    .Y(\soc/cpu/_01750_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_05997_  (.A1(\soc/cpu/_00711_ ),
    .A2(\soc/cpu/_01749_ ),
    .B1(\soc/cpu/_01750_ ),
    .Y(\soc/cpu/mem_la_addr [31]));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_05998_  (.A(\soc/cpu/is_compare ),
    .Y(\soc/cpu/_01751_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_05999_  (.A(\soc/cpu/instr_or ),
    .B(\soc/cpu/instr_ori ),
    .X(\soc/cpu/_01752_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06002_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/mem_la_wdata [0]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01755_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_06003_  (.A(\soc/cpu/instr_and ),
    .B(\soc/cpu/instr_andi ),
    .X(\soc/cpu/_01756_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_06006_  (.A(\soc/cpu/instr_xor ),
    .B(\soc/cpu/instr_xori ),
    .Y(\soc/cpu/_01759_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_06007_  (.A(\soc/cpu/instr_xor ),
    .B(\soc/cpu/instr_xori ),
    .X(\soc/cpu/_01760_ ));
 sky130_fd_sc_hd__or4_4 \soc/cpu/_06009_  (.A(\soc/cpu/is_compare ),
    .B(\soc/cpu/_01760_ ),
    .C(\soc/cpu/_01752_ ),
    .D(\soc/cpu/_01756_ ),
    .X(\soc/cpu/_01762_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06010_  (.A1(\soc/cpu/_01759_ ),
    .A2(\soc/cpu/_01762_ ),
    .B1(\soc/cpu/_01494_ ),
    .Y(\soc/cpu/_01763_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06011_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/mem_la_wdata [0]),
    .A3(\soc/cpu/_01756_ ),
    .B1(\soc/cpu/_01763_ ),
    .Y(\soc/cpu/_01764_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06012_  (.A1(\soc/cpu/_01751_ ),
    .A2(\soc/cpu/_01587_ ),
    .B1(\soc/cpu/_01755_ ),
    .C1(\soc/cpu/_01764_ ),
    .Y(\soc/cpu/alu_out[0] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06015_  (.A(\soc/cpu/mem_la_wdata [0]),
    .B(\soc/cpu/mem_la_wdata [1]),
    .Y(\soc/cpu/_01767_ ));
 sky130_fd_sc_hd__o21ba_1 \soc/cpu/_06016_  (.A1(\soc/cpu/mem_la_wdata [0]),
    .A2(\soc/cpu/mem_la_wdata [1]),
    .B1_N(\soc/cpu/instr_sub ),
    .X(\soc/cpu/_01768_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06017_  (.A1(\soc/cpu/instr_sub ),
    .A2(\soc/cpu/mem_la_wdata [1]),
    .B1(\soc/cpu/_01767_ ),
    .B2(\soc/cpu/_01768_ ),
    .Y(\soc/cpu/_01769_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06018_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/_01769_ ),
    .Y(\soc/cpu/_01770_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06019_  (.A(\soc/cpu/_01493_ ),
    .B(\soc/cpu/_01770_ ),
    .X(\soc/cpu/_01771_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06020_  (.A1(\soc/cpu/pcpi_rs1 [1]),
    .A2(net848),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01772_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06021_  (.A1(\soc/cpu/_01500_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01772_ ),
    .Y(\soc/cpu/_01773_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06022_  (.A1(net851),
    .A2(net848),
    .A3(\soc/cpu/_01756_ ),
    .B1(\soc/cpu/_01773_ ),
    .Y(\soc/cpu/_01774_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06023_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01771_ ),
    .B1(\soc/cpu/_01774_ ),
    .Y(\soc/cpu/alu_out[1] ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_06024_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/_01493_ ),
    .C(\soc/cpu/_01769_ ),
    .X(\soc/cpu/_01775_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06025_  (.A(\soc/cpu/mem_la_wdata [2]),
    .B(\soc/cpu/_01768_ ),
    .Y(\soc/cpu/_01776_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06026_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/_01776_ ),
    .X(\soc/cpu/_01777_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06027_  (.A(\soc/cpu/_01775_ ),
    .B(\soc/cpu/_01777_ ),
    .Y(\soc/cpu/_01778_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06028_  (.A1(\soc/cpu/pcpi_rs1 [2]),
    .A2(\soc/cpu/mem_la_wdata [2]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01779_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06030_  (.A1(\soc/cpu/_01507_ ),
    .A2(\soc/cpu/_01760_ ),
    .B1(\soc/cpu/_01756_ ),
    .B2(\soc/cpu/_01506_ ),
    .Y(\soc/cpu/_01781_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06031_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01778_ ),
    .B1(\soc/cpu/_01779_ ),
    .C1(\soc/cpu/_01781_ ),
    .Y(\soc/cpu/alu_out[2] ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_06032_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/_01775_ ),
    .C(\soc/cpu/_01776_ ),
    .X(\soc/cpu/_01782_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06033_  (.A(\soc/cpu/mem_la_wdata [0]),
    .B(\soc/cpu/mem_la_wdata [1]),
    .C(\soc/cpu/mem_la_wdata [2]),
    .Y(\soc/cpu/_01783_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06034_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01783_ ),
    .Y(\soc/cpu/_01784_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06035_  (.A(\soc/cpu/mem_la_wdata [3]),
    .B(\soc/cpu/_01784_ ),
    .Y(\soc/cpu/_01785_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06036_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(\soc/cpu/_01785_ ),
    .X(\soc/cpu/_01786_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06037_  (.A1(\soc/cpu/_01782_ ),
    .A2(\soc/cpu/_01786_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01787_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06038_  (.A1(\soc/cpu/_01782_ ),
    .A2(\soc/cpu/_01786_ ),
    .B1(\soc/cpu/_01787_ ),
    .Y(\soc/cpu/_01788_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06039_  (.A(\soc/cpu/_01503_ ),
    .B(\soc/cpu/_01760_ ),
    .Y(\soc/cpu/_01789_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06040_  (.A(net967),
    .B(\soc/cpu/mem_la_wdata [3]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01790_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06042_  (.A1(\soc/cpu/pcpi_rs1 [3]),
    .A2(\soc/cpu/mem_la_wdata [3]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01792_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_06043_  (.A(\soc/cpu/_01788_ ),
    .B(\soc/cpu/_01789_ ),
    .C(\soc/cpu/_01790_ ),
    .D(\soc/cpu/_01792_ ),
    .Y(\soc/cpu/alu_out[3] ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_06045_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(\soc/cpu/_01782_ ),
    .C(\soc/cpu/_01785_ ),
    .X(\soc/cpu/_01794_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06046_  (.A1(\soc/cpu/_01519_ ),
    .A2(\soc/cpu/_01783_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01795_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06047_  (.A(\soc/cpu/mem_la_wdata [4]),
    .B(\soc/cpu/_01795_ ),
    .Y(\soc/cpu/_01796_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06048_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/_01796_ ),
    .X(\soc/cpu/_01797_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06050_  (.A1(\soc/cpu/_01794_ ),
    .A2(\soc/cpu/_01797_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01799_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06051_  (.A1(\soc/cpu/_01794_ ),
    .A2(\soc/cpu/_01797_ ),
    .B1(\soc/cpu/_01799_ ),
    .Y(\soc/cpu/_01800_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06053_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/mem_la_wdata [4]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01802_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06055_  (.A1(\soc/cpu/pcpi_rs1 [4]),
    .A2(\soc/cpu/mem_la_wdata [4]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01804_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06056_  (.A1(\soc/cpu/_01498_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01800_ ),
    .C1(\soc/cpu/_01802_ ),
    .D1(\soc/cpu/_01804_ ),
    .Y(\soc/cpu/alu_out[4] ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_06057_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/_01794_ ),
    .C(\soc/cpu/_01796_ ),
    .X(\soc/cpu/_01805_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06058_  (.A(\soc/cpu/_01519_ ),
    .B(\soc/cpu/_01783_ ),
    .Y(\soc/cpu/_01806_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06059_  (.A(\soc/cpu/mem_la_wdata [4]),
    .B(\soc/cpu/_01806_ ),
    .Y(\soc/cpu/_01807_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06060_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01807_ ),
    .Y(\soc/cpu/_01808_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06061_  (.A(\soc/cpu/mem_la_wdata [5]),
    .B(\soc/cpu/_01808_ ),
    .Y(\soc/cpu/_01809_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06062_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(\soc/cpu/_01809_ ),
    .X(\soc/cpu/_01810_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06063_  (.A1(\soc/cpu/_01805_ ),
    .A2(\soc/cpu/_01810_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01811_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06064_  (.A1(\soc/cpu/_01805_ ),
    .A2(\soc/cpu/_01810_ ),
    .B1(\soc/cpu/_01811_ ),
    .Y(\soc/cpu/_01812_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06065_  (.A(net860),
    .B(\soc/cpu/mem_la_wdata [5]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01813_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06066_  (.A1(net860),
    .A2(\soc/cpu/mem_la_wdata [5]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01814_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06067_  (.A1(\soc/cpu/_01496_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01812_ ),
    .C1(\soc/cpu/_01813_ ),
    .D1(\soc/cpu/_01814_ ),
    .Y(\soc/cpu/alu_out[5] ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_06068_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(\soc/cpu/_01805_ ),
    .C(\soc/cpu/_01809_ ),
    .X(\soc/cpu/_01815_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06069_  (.A1(\soc/cpu/_01517_ ),
    .A2(\soc/cpu/_01807_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01816_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06070_  (.A(net788),
    .B(\soc/cpu/_01816_ ),
    .Y(\soc/cpu/_01817_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06071_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(\soc/cpu/_01817_ ),
    .X(\soc/cpu/_01818_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06072_  (.A1(\soc/cpu/_01815_ ),
    .A2(\soc/cpu/_01818_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01819_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06073_  (.A1(\soc/cpu/_01815_ ),
    .A2(\soc/cpu/_01818_ ),
    .B1(\soc/cpu/_01819_ ),
    .Y(\soc/cpu/_01820_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06074_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(net776),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01821_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06075_  (.A1(\soc/cpu/pcpi_rs1 [6]),
    .A2(net776),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01822_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06076_  (.A1(\soc/cpu/_01510_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01820_ ),
    .C1(\soc/cpu/_01821_ ),
    .D1(\soc/cpu/_01822_ ),
    .Y(\soc/cpu/alu_out[6] ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_06077_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(\soc/cpu/_01815_ ),
    .C(\soc/cpu/_01817_ ),
    .X(\soc/cpu/_01823_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_06078_  (.A(\soc/cpu/mem_la_wdata [5]),
    .B(\soc/cpu/mem_la_wdata [4]),
    .C(\soc/cpu/mem_la_wdata [6]),
    .D(\soc/cpu/_01806_ ),
    .Y(\soc/cpu/_01824_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06079_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01824_ ),
    .Y(\soc/cpu/_01825_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06080_  (.A(net773),
    .B(\soc/cpu/_01825_ ),
    .Y(\soc/cpu/_01826_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06081_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(\soc/cpu/_01826_ ),
    .X(\soc/cpu/_01827_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06082_  (.A(\soc/cpu/_01823_ ),
    .B(\soc/cpu/_01827_ ),
    .Y(\soc/cpu/_01828_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06083_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(net773),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01829_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06085_  (.A1(\soc/cpu/pcpi_rs1 [7]),
    .A2(net773),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01831_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06086_  (.A1(\soc/cpu/pcpi_rs1 [7]),
    .A2(net773),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01831_ ),
    .Y(\soc/cpu/_01832_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06087_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01828_ ),
    .B1(net774),
    .C1(\soc/cpu/_01832_ ),
    .Y(\soc/cpu/alu_out[7] ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06088_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(net780),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01833_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06089_  (.A1(\soc/cpu/pcpi_rs1 [8]),
    .A2(net780),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01834_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06090_  (.A1(\soc/cpu/pcpi_rs1 [8]),
    .A2(net780),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01834_ ),
    .Y(\soc/cpu/_01835_ ));
 sky130_fd_sc_hd__maj3_2 \soc/cpu/_06091_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(\soc/cpu/_01823_ ),
    .C(\soc/cpu/_01826_ ),
    .X(\soc/cpu/_01836_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06092_  (.A1(\soc/cpu/_01516_ ),
    .A2(\soc/cpu/_01824_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01837_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06093_  (.A(\soc/cpu/pcpi_rs2 [8]),
    .B(\soc/cpu/_01837_ ),
    .Y(\soc/cpu/_01838_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06094_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(\soc/cpu/_01838_ ),
    .X(\soc/cpu/_01839_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06095_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(\soc/cpu/_01838_ ),
    .Y(\soc/cpu/_01840_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06096_  (.A(\soc/cpu/_01839_ ),
    .B(\soc/cpu/_01840_ ),
    .Y(\soc/cpu/_01841_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06097_  (.A1(\soc/cpu/_01836_ ),
    .A2(\soc/cpu/_01841_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01842_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06098_  (.A1(\soc/cpu/_01836_ ),
    .A2(\soc/cpu/_01841_ ),
    .B1(\soc/cpu/_01842_ ),
    .Y(\soc/cpu/_01843_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06099_  (.A(\soc/cpu/_01833_ ),
    .B(\soc/cpu/_01835_ ),
    .C(\soc/cpu/_01843_ ),
    .Y(\soc/cpu/alu_out[8] ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_06100_  (.A1(\soc/cpu/_01836_ ),
    .A2(\soc/cpu/_01841_ ),
    .B1(\soc/cpu/_01839_ ),
    .X(\soc/cpu/_01844_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06101_  (.A(net780),
    .Y(\soc/cpu/_01845_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06102_  (.A1(\soc/cpu/_01516_ ),
    .A2(\soc/cpu/_01845_ ),
    .A3(\soc/cpu/_01824_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01846_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06103_  (.A(\soc/cpu/pcpi_rs2 [9]),
    .B(\soc/cpu/_01846_ ),
    .Y(\soc/cpu/_01847_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06104_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(\soc/cpu/_01847_ ),
    .X(\soc/cpu/_01848_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06105_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(\soc/cpu/_01847_ ),
    .Y(\soc/cpu/_01849_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06106_  (.A(\soc/cpu/_01848_ ),
    .B(\soc/cpu/_01849_ ),
    .Y(\soc/cpu/_01850_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06107_  (.A1(\soc/cpu/_01844_ ),
    .A2(\soc/cpu/_01850_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01851_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06108_  (.A1(\soc/cpu/_01844_ ),
    .A2(\soc/cpu/_01850_ ),
    .B1(\soc/cpu/_01851_ ),
    .Y(\soc/cpu/_01852_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06109_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(net781),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01853_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06110_  (.A1(\soc/cpu/pcpi_rs1 [9]),
    .A2(net781),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01854_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06111_  (.A1(\soc/cpu/_01475_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01852_ ),
    .C1(\soc/cpu/_01853_ ),
    .D1(\soc/cpu/_01854_ ),
    .Y(\soc/cpu/alu_out[9] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06112_  (.A(\soc/cpu/_01516_ ),
    .B(\soc/cpu/_01824_ ),
    .Y(\soc/cpu/_01855_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_06113_  (.A(\soc/cpu/pcpi_rs2 [9]),
    .B(\soc/cpu/pcpi_rs2 [8]),
    .C(\soc/cpu/_01855_ ),
    .Y(\soc/cpu/_01856_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06114_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01856_ ),
    .Y(\soc/cpu/_01857_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06115_  (.A(\soc/cpu/pcpi_rs2 [10]),
    .B(\soc/cpu/_01857_ ),
    .Y(\soc/cpu/_01858_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06116_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(\soc/cpu/_01858_ ),
    .Y(\soc/cpu/_01859_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06117_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(\soc/cpu/_01858_ ),
    .Y(\soc/cpu/_01860_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_06118_  (.A(\soc/cpu/_01859_ ),
    .SLEEP(\soc/cpu/_01860_ ),
    .X(\soc/cpu/_01861_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_06119_  (.A1(\soc/cpu/_01836_ ),
    .A2(\soc/cpu/_01841_ ),
    .B1(\soc/cpu/_01848_ ),
    .C1(\soc/cpu/_01839_ ),
    .Y(\soc/cpu/_01862_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06120_  (.A(\soc/cpu/_01849_ ),
    .B(\soc/cpu/_01862_ ),
    .Y(\soc/cpu/_01863_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06121_  (.A(\soc/cpu/_01861_ ),
    .B(\soc/cpu/_01863_ ),
    .Y(\soc/cpu/_01864_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06122_  (.A1(\soc/cpu/pcpi_rs1 [10]),
    .A2(\soc/cpu/pcpi_rs2 [10]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01865_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06123_  (.A1(\soc/cpu/pcpi_rs1 [10]),
    .A2(\soc/cpu/pcpi_rs2 [10]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01865_ ),
    .Y(\soc/cpu/_01866_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06124_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(\soc/cpu/pcpi_rs2 [10]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01867_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06125_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01864_ ),
    .B1(\soc/cpu/_01866_ ),
    .C1(\soc/cpu/_01867_ ),
    .Y(\soc/cpu/alu_out[10] ));
 sky130_fd_sc_hd__o31ai_2 \soc/cpu/_06126_  (.A1(\soc/cpu/_01849_ ),
    .A2(\soc/cpu/_01860_ ),
    .A3(\soc/cpu/_01862_ ),
    .B1(\soc/cpu/_01859_ ),
    .Y(\soc/cpu/_01868_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_06127_  (.A(\soc/cpu/pcpi_rs2 [10]),
    .Y(\soc/cpu/_01869_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06128_  (.A1(\soc/cpu/_01869_ ),
    .A2(\soc/cpu/_01856_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01870_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06129_  (.A(net777),
    .B(\soc/cpu/_01870_ ),
    .Y(\soc/cpu/_01871_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06130_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(\soc/cpu/_01871_ ),
    .X(\soc/cpu/_01872_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06131_  (.A(\soc/cpu/_01868_ ),
    .B(\soc/cpu/_01872_ ),
    .Y(\soc/cpu/_01873_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06132_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(net777),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01874_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06133_  (.A1(\soc/cpu/pcpi_rs1 [11]),
    .A2(net777),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01875_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06134_  (.A1(\soc/cpu/pcpi_rs1 [11]),
    .A2(net777),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01875_ ),
    .Y(\soc/cpu/_01876_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06135_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01873_ ),
    .B1(\soc/cpu/_01874_ ),
    .C1(\soc/cpu/_01876_ ),
    .Y(\soc/cpu/alu_out[11] ));
 sky130_fd_sc_hd__maj3_2 \soc/cpu/_06136_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(\soc/cpu/_01868_ ),
    .C(\soc/cpu/_01871_ ),
    .X(\soc/cpu/_01877_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06137_  (.A1(\soc/cpu/_01537_ ),
    .A2(\soc/cpu/_01869_ ),
    .A3(\soc/cpu/_01856_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01878_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06138_  (.A(\soc/cpu/pcpi_rs2 [12]),
    .B(\soc/cpu/_01878_ ),
    .Y(\soc/cpu/_01879_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06139_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/_01879_ ),
    .X(\soc/cpu/_01880_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06140_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/_01879_ ),
    .Y(\soc/cpu/_01881_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06141_  (.A(\soc/cpu/_01880_ ),
    .B(\soc/cpu/_01881_ ),
    .Y(\soc/cpu/_01882_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06142_  (.A(\soc/cpu/_01877_ ),
    .B(\soc/cpu/_01882_ ),
    .Y(\soc/cpu/_01883_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06143_  (.A1(\soc/cpu/pcpi_rs1 [12]),
    .A2(\soc/cpu/pcpi_rs2 [12]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01884_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06144_  (.A1(\soc/cpu/pcpi_rs1 [12]),
    .A2(\soc/cpu/pcpi_rs2 [12]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01884_ ),
    .Y(\soc/cpu/_01885_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06145_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/pcpi_rs2 [12]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01886_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06146_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01883_ ),
    .B1(\soc/cpu/_01885_ ),
    .C1(\soc/cpu/_01886_ ),
    .Y(\soc/cpu/alu_out[12] ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06147_  (.A(\soc/cpu/_01877_ ),
    .B(\soc/cpu/_01882_ ),
    .X(\soc/cpu/_01887_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06148_  (.A(\soc/cpu/_01869_ ),
    .B(\soc/cpu/_01856_ ),
    .Y(\soc/cpu/_01888_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_06149_  (.A(\soc/cpu/pcpi_rs2 [11]),
    .B(\soc/cpu/pcpi_rs2 [12]),
    .C(\soc/cpu/_01888_ ),
    .Y(\soc/cpu/_01889_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06150_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01889_ ),
    .Y(\soc/cpu/_01890_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06151_  (.A(\soc/cpu/pcpi_rs2 [13]),
    .B(\soc/cpu/_01890_ ),
    .Y(\soc/cpu/_01891_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06152_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/_01891_ ),
    .X(\soc/cpu/_01892_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06153_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/_01891_ ),
    .Y(\soc/cpu/_01893_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06154_  (.A(\soc/cpu/_01892_ ),
    .B(\soc/cpu/_01893_ ),
    .Y(\soc/cpu/_01894_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_06155_  (.A1(\soc/cpu/_01880_ ),
    .A2(\soc/cpu/_01887_ ),
    .B1(\soc/cpu/_01894_ ),
    .X(\soc/cpu/_01895_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_06156_  (.A(\soc/cpu/is_compare ),
    .B(\soc/cpu/_01760_ ),
    .C(\soc/cpu/_01752_ ),
    .D(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01896_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06157_  (.A1(\soc/cpu/_01880_ ),
    .A2(\soc/cpu/_01887_ ),
    .A3(\soc/cpu/_01894_ ),
    .B1(net145),
    .Y(\soc/cpu/_01897_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06158_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/pcpi_rs2 [13]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01898_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06159_  (.A1(\soc/cpu/pcpi_rs1 [13]),
    .A2(\soc/cpu/pcpi_rs2 [13]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01899_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06160_  (.A1(\soc/cpu/pcpi_rs1 [13]),
    .A2(\soc/cpu/pcpi_rs2 [13]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01899_ ),
    .Y(\soc/cpu/_01900_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06161_  (.A1(\soc/cpu/_01895_ ),
    .A2(\soc/cpu/_01897_ ),
    .B1(\soc/cpu/_01898_ ),
    .C1(\soc/cpu/_01900_ ),
    .Y(\soc/cpu/alu_out[13] ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_06162_  (.A1(\soc/cpu/_01877_ ),
    .A2(\soc/cpu/_01882_ ),
    .B1(\soc/cpu/_01892_ ),
    .C1(\soc/cpu/_01880_ ),
    .Y(\soc/cpu/_01901_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06163_  (.A1(\soc/cpu/_01533_ ),
    .A2(\soc/cpu/_01889_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01902_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06164_  (.A(\soc/cpu/pcpi_rs2 [14]),
    .B(\soc/cpu/_01902_ ),
    .Y(\soc/cpu/_01903_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06165_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(\soc/cpu/_01903_ ),
    .Y(\soc/cpu/_01904_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_06166_  (.A1(\soc/cpu/_01893_ ),
    .A2(\soc/cpu/_01901_ ),
    .B1(\soc/cpu/_01904_ ),
    .X(\soc/cpu/_01905_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06167_  (.A1(\soc/cpu/_01893_ ),
    .A2(\soc/cpu/_01904_ ),
    .A3(\soc/cpu/_01901_ ),
    .B1(net145),
    .Y(\soc/cpu/_01906_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06168_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(\soc/cpu/pcpi_rs2 [14]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01907_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06169_  (.A1(\soc/cpu/pcpi_rs1 [14]),
    .A2(\soc/cpu/pcpi_rs2 [14]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01908_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06170_  (.A1(\soc/cpu/pcpi_rs1 [14]),
    .A2(\soc/cpu/pcpi_rs2 [14]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01908_ ),
    .Y(\soc/cpu/_01909_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06171_  (.A1(\soc/cpu/_01905_ ),
    .A2(\soc/cpu/_01906_ ),
    .B1(\soc/cpu/_01907_ ),
    .C1(\soc/cpu/_01909_ ),
    .Y(\soc/cpu/alu_out[14] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06172_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(\soc/cpu/_01903_ ),
    .Y(\soc/cpu/_01910_ ));
 sky130_fd_sc_hd__o31ai_2 \soc/cpu/_06173_  (.A1(\soc/cpu/_01893_ ),
    .A2(\soc/cpu/_01904_ ),
    .A3(\soc/cpu/_01901_ ),
    .B1(\soc/cpu/_01910_ ),
    .Y(\soc/cpu/_01911_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06174_  (.A(\soc/cpu/pcpi_rs2 [14]),
    .Y(\soc/cpu/_01912_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06175_  (.A1(\soc/cpu/_01533_ ),
    .A2(\soc/cpu/_01912_ ),
    .A3(\soc/cpu/_01889_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01913_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06176_  (.A(\soc/cpu/pcpi_rs2 [15]),
    .B(\soc/cpu/_01913_ ),
    .Y(\soc/cpu/_01914_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06177_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(\soc/cpu/_01914_ ),
    .X(\soc/cpu/_01915_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06178_  (.A1(\soc/cpu/_01911_ ),
    .A2(\soc/cpu/_01915_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01916_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06179_  (.A1(\soc/cpu/_01911_ ),
    .A2(\soc/cpu/_01915_ ),
    .B1(\soc/cpu/_01916_ ),
    .Y(\soc/cpu/_01917_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06180_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(\soc/cpu/pcpi_rs2 [15]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01918_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06181_  (.A1(\soc/cpu/pcpi_rs1 [15]),
    .A2(\soc/cpu/pcpi_rs2 [15]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01919_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06182_  (.A1(\soc/cpu/_01478_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01917_ ),
    .C1(\soc/cpu/_01918_ ),
    .D1(\soc/cpu/_01919_ ),
    .Y(\soc/cpu/alu_out[15] ));
 sky130_fd_sc_hd__maj3_2 \soc/cpu/_06183_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(\soc/cpu/_01911_ ),
    .C(\soc/cpu/_01914_ ),
    .X(\soc/cpu/_01920_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06184_  (.A(\soc/cpu/_01533_ ),
    .B(\soc/cpu/_01889_ ),
    .Y(\soc/cpu/_01921_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06185_  (.A(\soc/cpu/pcpi_rs2 [15]),
    .B(\soc/cpu/pcpi_rs2 [14]),
    .C(\soc/cpu/_01921_ ),
    .Y(\soc/cpu/_01922_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06186_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01922_ ),
    .Y(\soc/cpu/_01923_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06187_  (.A(\soc/cpu/pcpi_rs2 [16]),
    .B(\soc/cpu/_01923_ ),
    .Y(\soc/cpu/_01924_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06188_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(\soc/cpu/_01924_ ),
    .X(\soc/cpu/_01925_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06189_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(\soc/cpu/_01924_ ),
    .Y(\soc/cpu/_01926_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06190_  (.A(\soc/cpu/_01925_ ),
    .B(\soc/cpu/_01926_ ),
    .Y(\soc/cpu/_01927_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06191_  (.A(\soc/cpu/_01920_ ),
    .B(\soc/cpu/_01927_ ),
    .Y(\soc/cpu/_01928_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06192_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(\soc/cpu/pcpi_rs2 [16]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01929_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06193_  (.A1(\soc/cpu/pcpi_rs1 [16]),
    .A2(\soc/cpu/pcpi_rs2 [16]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01930_ ));
 sky130_fd_sc_hd__o211a_1 \soc/cpu/_06194_  (.A1(\soc/cpu/_01453_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01929_ ),
    .C1(\soc/cpu/_01930_ ),
    .X(\soc/cpu/_01931_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06195_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01928_ ),
    .B1(\soc/cpu/_01931_ ),
    .Y(\soc/cpu/alu_out[16] ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_06196_  (.A1(\soc/cpu/_01920_ ),
    .A2(\soc/cpu/_01927_ ),
    .B1(\soc/cpu/_01925_ ),
    .X(\soc/cpu/_01932_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06197_  (.A_N(\soc/cpu/pcpi_rs2 [16]),
    .B(\soc/cpu/_01922_ ),
    .Y(\soc/cpu/_01933_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_06198_  (.A(\soc/cpu/instr_sub ),
    .B_N(\soc/cpu/_01933_ ),
    .Y(\soc/cpu/_01934_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06199_  (.A(\soc/cpu/pcpi_rs2 [17]),
    .B(\soc/cpu/_01934_ ),
    .Y(\soc/cpu/_01935_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06200_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(\soc/cpu/_01935_ ),
    .X(\soc/cpu/_01936_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06201_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(\soc/cpu/_01935_ ),
    .Y(\soc/cpu/_01937_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06202_  (.A(\soc/cpu/_01936_ ),
    .B(\soc/cpu/_01937_ ),
    .Y(\soc/cpu/_01938_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06203_  (.A1(\soc/cpu/_01932_ ),
    .A2(\soc/cpu/_01938_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_01939_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06204_  (.A1(\soc/cpu/_01932_ ),
    .A2(\soc/cpu/_01938_ ),
    .B1(\soc/cpu/_01939_ ),
    .Y(\soc/cpu/_01940_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06205_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(\soc/cpu/pcpi_rs2 [17]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01941_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06206_  (.A1(\soc/cpu/pcpi_rs1 [17]),
    .A2(\soc/cpu/pcpi_rs2 [17]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01942_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06207_  (.A1(\soc/cpu/_01448_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01940_ ),
    .C1(\soc/cpu/_01941_ ),
    .D1(\soc/cpu/_01942_ ),
    .Y(\soc/cpu/alu_out[17] ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06208_  (.A(\soc/cpu/pcpi_rs2 [17]),
    .B(\soc/cpu/_01933_ ),
    .Y(\soc/cpu/_01943_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06209_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01943_ ),
    .Y(\soc/cpu/_01944_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06210_  (.A(\soc/cpu/pcpi_rs2 [18]),
    .B(\soc/cpu/_01944_ ),
    .Y(\soc/cpu/_01945_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06211_  (.A(\soc/cpu/_01555_ ),
    .B(\soc/cpu/_01945_ ),
    .Y(\soc/cpu/_01946_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/cpu/_06212_  (.A1(\soc/cpu/_01920_ ),
    .A2(\soc/cpu/_01927_ ),
    .B1(\soc/cpu/_01936_ ),
    .C1(\soc/cpu/_01925_ ),
    .Y(\soc/cpu/_01947_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06213_  (.A(\soc/cpu/_01937_ ),
    .B(\soc/cpu/_01947_ ),
    .Y(\soc/cpu/_01948_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06214_  (.A(\soc/cpu/_01946_ ),
    .B(\soc/cpu/_01948_ ),
    .Y(\soc/cpu/_01949_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06215_  (.A(\soc/cpu/pcpi_rs1 [18]),
    .B(\soc/cpu/pcpi_rs2 [18]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01950_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06216_  (.A1(\soc/cpu/pcpi_rs1 [18]),
    .A2(\soc/cpu/pcpi_rs2 [18]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01951_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06217_  (.A1(\soc/cpu/pcpi_rs1 [18]),
    .A2(\soc/cpu/pcpi_rs2 [18]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01951_ ),
    .Y(\soc/cpu/_01952_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06218_  (.A1(\soc/cpu/_01762_ ),
    .A2(\soc/cpu/_01949_ ),
    .B1(\soc/cpu/_01950_ ),
    .C1(\soc/cpu/_01952_ ),
    .Y(\soc/cpu/alu_out[18] ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06219_  (.A(\soc/cpu/_01946_ ),
    .Y(\soc/cpu/_01953_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06220_  (.A(\soc/cpu/pcpi_rs1 [18]),
    .B(\soc/cpu/_01945_ ),
    .Y(\soc/cpu/_01954_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06221_  (.A1(\soc/cpu/_01937_ ),
    .A2(\soc/cpu/_01953_ ),
    .A3(\soc/cpu/_01947_ ),
    .B1(\soc/cpu/_01954_ ),
    .Y(\soc/cpu/_01955_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06222_  (.A(\soc/cpu/pcpi_rs2 [18]),
    .B(\soc/cpu/pcpi_rs2 [17]),
    .C(\soc/cpu/_01933_ ),
    .Y(\soc/cpu/_01956_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06223_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01956_ ),
    .Y(\soc/cpu/_01957_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06224_  (.A(\soc/cpu/pcpi_rs2 [19]),
    .B(\soc/cpu/_01957_ ),
    .Y(\soc/cpu/_01958_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06225_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(\soc/cpu/_01958_ ),
    .Y(\soc/cpu/_01959_ ));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_06226_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(\soc/cpu/_01958_ ),
    .X(\soc/cpu/_01960_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06227_  (.A(\soc/cpu/_01959_ ),
    .B(\soc/cpu/_01960_ ),
    .Y(\soc/cpu/_01961_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06228_  (.A(\soc/cpu/_01955_ ),
    .B(\soc/cpu/_01961_ ),
    .Y(\soc/cpu/_01962_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06229_  (.A(net145),
    .B(\soc/cpu/_01962_ ),
    .Y(\soc/cpu/_01963_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06230_  (.A(net881),
    .B(\soc/cpu/pcpi_rs2 [19]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01964_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06231_  (.A1(\soc/cpu/pcpi_rs1 [19]),
    .A2(\soc/cpu/pcpi_rs2 [19]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01965_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06232_  (.A1(\soc/cpu/_01454_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01963_ ),
    .C1(\soc/cpu/_01964_ ),
    .D1(\soc/cpu/_01965_ ),
    .Y(\soc/cpu/alu_out[19] ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06233_  (.A(\soc/cpu/pcpi_rs1 [20]),
    .B(\soc/cpu/pcpi_rs2 [20]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01966_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06234_  (.A1(\soc/cpu/pcpi_rs1 [20]),
    .A2(\soc/cpu/pcpi_rs2 [20]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01967_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06235_  (.A1(\soc/cpu/pcpi_rs1 [20]),
    .A2(\soc/cpu/pcpi_rs2 [20]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01967_ ),
    .Y(\soc/cpu/_01968_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06236_  (.A1(\soc/cpu/_01554_ ),
    .A2(\soc/cpu/_01956_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_01969_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06237_  (.A(\soc/cpu/pcpi_rs2 [20]),
    .B(\soc/cpu/_01969_ ),
    .Y(\soc/cpu/_01970_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06238_  (.A(\soc/cpu/pcpi_rs1 [20]),
    .B(\soc/cpu/_01970_ ),
    .X(\soc/cpu/_01971_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06239_  (.A(\soc/cpu/pcpi_rs1 [20]),
    .B(\soc/cpu/_01970_ ),
    .Y(\soc/cpu/_01972_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06240_  (.A(\soc/cpu/_01971_ ),
    .B(\soc/cpu/_01972_ ),
    .Y(\soc/cpu/_01973_ ));
 sky130_fd_sc_hd__o311ai_4 \soc/cpu/_06241_  (.A1(\soc/cpu/_01937_ ),
    .A2(\soc/cpu/_01953_ ),
    .A3(\soc/cpu/_01947_ ),
    .B1(\soc/cpu/_01959_ ),
    .C1(\soc/cpu/_01954_ ),
    .Y(\soc/cpu/_01974_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06242_  (.A1(\soc/cpu/_01960_ ),
    .A2(\soc/cpu/_01974_ ),
    .B1(\soc/cpu/_01973_ ),
    .Y(\soc/cpu/_01975_ ));
 sky130_fd_sc_hd__a311o_1 \soc/cpu/_06243_  (.A1(\soc/cpu/_01960_ ),
    .A2(\soc/cpu/_01973_ ),
    .A3(\soc/cpu/_01974_ ),
    .B1(\soc/cpu/_01975_ ),
    .C1(\soc/cpu/_01762_ ),
    .X(\soc/cpu/_01976_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06244_  (.A(\soc/cpu/_01966_ ),
    .B(\soc/cpu/_01968_ ),
    .C(\soc/cpu/_01976_ ),
    .Y(\soc/cpu/alu_out[20] ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06245_  (.A1(\soc/cpu/_01960_ ),
    .A2(\soc/cpu/_01973_ ),
    .A3(\soc/cpu/_01974_ ),
    .B1(\soc/cpu/_01971_ ),
    .Y(\soc/cpu/_01977_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06246_  (.A(\soc/cpu/_01554_ ),
    .B(\soc/cpu/_01956_ ),
    .Y(\soc/cpu/_01978_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06247_  (.A(\soc/cpu/pcpi_rs2 [20]),
    .B(\soc/cpu/_01978_ ),
    .Y(\soc/cpu/_01979_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06248_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01979_ ),
    .Y(\soc/cpu/_01980_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06249_  (.A(\soc/cpu/pcpi_rs2 [21]),
    .B(\soc/cpu/_01980_ ),
    .Y(\soc/cpu/_01981_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06250_  (.A(\soc/cpu/pcpi_rs1 [21]),
    .B(\soc/cpu/_01981_ ),
    .X(\soc/cpu/_01982_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06251_  (.A(\soc/cpu/pcpi_rs1 [21]),
    .B(\soc/cpu/_01981_ ),
    .Y(\soc/cpu/_01983_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06252_  (.A(\soc/cpu/_01982_ ),
    .B(\soc/cpu/_01983_ ),
    .Y(\soc/cpu/_01984_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06253_  (.A(\soc/cpu/_01977_ ),
    .B(\soc/cpu/_01984_ ),
    .Y(\soc/cpu/_01985_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06254_  (.A(net145),
    .B(\soc/cpu/_01985_ ),
    .Y(\soc/cpu/_01986_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06255_  (.A(net893),
    .B(\soc/cpu/pcpi_rs2 [21]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01987_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06256_  (.A1(\soc/cpu/pcpi_rs1 [21]),
    .A2(\soc/cpu/pcpi_rs2 [21]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_01988_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06257_  (.A1(\soc/cpu/_01456_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_01986_ ),
    .C1(\soc/cpu/_01987_ ),
    .D1(\soc/cpu/_01988_ ),
    .Y(\soc/cpu/alu_out[21] ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06258_  (.A(\soc/cpu/pcpi_rs2 [21]),
    .B(\soc/cpu/pcpi_rs2 [20]),
    .C(\soc/cpu/_01978_ ),
    .Y(\soc/cpu/_01989_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06259_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_01989_ ),
    .Y(\soc/cpu/_01990_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_06260_  (.A(net754),
    .B(\soc/cpu/_01990_ ),
    .Y(\soc/cpu/_01991_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_06261_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(\soc/cpu/_01991_ ),
    .Y(\soc/cpu/_01992_ ));
 sky130_fd_sc_hd__a311oi_4 \soc/cpu/_06262_  (.A1(\soc/cpu/_01960_ ),
    .A2(\soc/cpu/_01973_ ),
    .A3(\soc/cpu/_01974_ ),
    .B1(\soc/cpu/_01982_ ),
    .C1(\soc/cpu/_01971_ ),
    .Y(\soc/cpu/_01993_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06263_  (.A(\soc/cpu/_01983_ ),
    .B(\soc/cpu/_01992_ ),
    .C(\soc/cpu/_01993_ ),
    .Y(\soc/cpu/_01994_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06264_  (.A1(\soc/cpu/_01983_ ),
    .A2(\soc/cpu/_01993_ ),
    .B1(\soc/cpu/_01992_ ),
    .Y(\soc/cpu/_01995_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06265_  (.A(net145),
    .B(\soc/cpu/_01995_ ),
    .Y(\soc/cpu/_01996_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06266_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(net754),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_01997_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06267_  (.A1(\soc/cpu/pcpi_rs1 [22]),
    .A2(net754),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_01998_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06268_  (.A1(\soc/cpu/pcpi_rs1 [22]),
    .A2(net754),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_01998_ ),
    .Y(\soc/cpu/_01999_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06269_  (.A1(\soc/cpu/_01994_ ),
    .A2(\soc/cpu/_01996_ ),
    .B1(net755),
    .C1(\soc/cpu/_01999_ ),
    .Y(\soc/cpu/alu_out[22] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06270_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(\soc/cpu/_01991_ ),
    .Y(\soc/cpu/_02000_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06271_  (.A1(\soc/cpu/_01983_ ),
    .A2(\soc/cpu/_01992_ ),
    .A3(\soc/cpu/_01993_ ),
    .B1(\soc/cpu/_02000_ ),
    .Y(\soc/cpu/_02001_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06272_  (.A_N(\soc/cpu/pcpi_rs2 [22]),
    .B(\soc/cpu/_01989_ ),
    .Y(\soc/cpu/_02002_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_06273_  (.A(\soc/cpu/instr_sub ),
    .B_N(\soc/cpu/_02002_ ),
    .Y(\soc/cpu/_02003_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06274_  (.A(\soc/cpu/pcpi_rs2 [23]),
    .B(\soc/cpu/_02003_ ),
    .Y(\soc/cpu/_02004_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06275_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(\soc/cpu/_02004_ ),
    .Y(\soc/cpu/_02005_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_06276_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(\soc/cpu/_02004_ ),
    .X(\soc/cpu/_02006_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06277_  (.A(\soc/cpu/_02005_ ),
    .B(\soc/cpu/_02006_ ),
    .X(\soc/cpu/_02007_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06278_  (.A1(\soc/cpu/_02001_ ),
    .A2(\soc/cpu/_02007_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_02008_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06279_  (.A1(\soc/cpu/_02001_ ),
    .A2(\soc/cpu/_02007_ ),
    .B1(\soc/cpu/_02008_ ),
    .Y(\soc/cpu/_02009_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06280_  (.A(net895),
    .B(\soc/cpu/pcpi_rs2 [23]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02010_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06281_  (.A1(\soc/cpu/pcpi_rs1 [23]),
    .A2(\soc/cpu/pcpi_rs2 [23]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_02011_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06282_  (.A1(\soc/cpu/_01458_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_02009_ ),
    .C1(\soc/cpu/_02010_ ),
    .D1(\soc/cpu/_02011_ ),
    .Y(\soc/cpu/alu_out[23] ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06283_  (.A(\soc/cpu/pcpi_rs2 [23]),
    .B(\soc/cpu/_02002_ ),
    .Y(\soc/cpu/_02012_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06284_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_02012_ ),
    .Y(\soc/cpu/_02013_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06285_  (.A(\soc/cpu/pcpi_rs2 [24]),
    .B(\soc/cpu/_02013_ ),
    .Y(\soc/cpu/_02014_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06286_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(\soc/cpu/_02014_ ),
    .X(\soc/cpu/_02015_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06287_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(\soc/cpu/_02014_ ),
    .Y(\soc/cpu/_02016_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06288_  (.A(\soc/cpu/_02015_ ),
    .B(\soc/cpu/_02016_ ),
    .Y(\soc/cpu/_02017_ ));
 sky130_fd_sc_hd__o311ai_4 \soc/cpu/_06289_  (.A1(\soc/cpu/_01983_ ),
    .A2(\soc/cpu/_01992_ ),
    .A3(\soc/cpu/_01993_ ),
    .B1(\soc/cpu/_02005_ ),
    .C1(\soc/cpu/_02000_ ),
    .Y(\soc/cpu/_02018_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06290_  (.A(\soc/cpu/_02006_ ),
    .B(\soc/cpu/_02018_ ),
    .X(\soc/cpu/_02019_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06291_  (.A1(\soc/cpu/_02017_ ),
    .A2(\soc/cpu/_02019_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_02020_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06292_  (.A1(\soc/cpu/_02017_ ),
    .A2(\soc/cpu/_02019_ ),
    .B1(\soc/cpu/_02020_ ),
    .Y(\soc/cpu/_02021_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06293_  (.A(\soc/cpu/_01439_ ),
    .B(\soc/cpu/_01760_ ),
    .Y(\soc/cpu/_02022_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06294_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(\soc/cpu/pcpi_rs2 [24]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02023_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06295_  (.A1(\soc/cpu/pcpi_rs1 [24]),
    .A2(\soc/cpu/pcpi_rs2 [24]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_02024_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_06296_  (.A(\soc/cpu/_02021_ ),
    .B(\soc/cpu/_02022_ ),
    .C(\soc/cpu/_02023_ ),
    .D(\soc/cpu/_02024_ ),
    .Y(\soc/cpu/alu_out[24] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06297_  (.A1(\soc/cpu/_02017_ ),
    .A2(\soc/cpu/_02019_ ),
    .B1(\soc/cpu/_02015_ ),
    .Y(\soc/cpu/_02025_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06298_  (.A(\soc/cpu/pcpi_rs2 [24]),
    .B(\soc/cpu/pcpi_rs2 [23]),
    .C(\soc/cpu/_02002_ ),
    .Y(\soc/cpu/_02026_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06299_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_02026_ ),
    .Y(\soc/cpu/_02027_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06300_  (.A(\soc/cpu/pcpi_rs2 [25]),
    .B(\soc/cpu/_02027_ ),
    .Y(\soc/cpu/_02028_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06301_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .B(\soc/cpu/_02028_ ),
    .X(\soc/cpu/_02029_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06302_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .B(\soc/cpu/_02028_ ),
    .Y(\soc/cpu/_02030_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06303_  (.A(\soc/cpu/_02029_ ),
    .B(\soc/cpu/_02030_ ),
    .Y(\soc/cpu/_02031_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06304_  (.A(\soc/cpu/_02025_ ),
    .B(\soc/cpu/_02031_ ),
    .Y(\soc/cpu/_02032_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06305_  (.A(net145),
    .B(\soc/cpu/_02032_ ),
    .Y(\soc/cpu/_02033_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06306_  (.A(\soc/cpu/_01433_ ),
    .B(\soc/cpu/_01760_ ),
    .Y(\soc/cpu/_02034_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06307_  (.A(net897),
    .B(\soc/cpu/pcpi_rs2 [25]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02035_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06308_  (.A1(\soc/cpu/pcpi_rs1 [25]),
    .A2(\soc/cpu/pcpi_rs2 [25]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_02036_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_06309_  (.A(\soc/cpu/_02033_ ),
    .B(\soc/cpu/_02034_ ),
    .C(\soc/cpu/_02035_ ),
    .D(\soc/cpu/_02036_ ),
    .Y(\soc/cpu/alu_out[25] ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06310_  (.A(\soc/cpu/pcpi_rs2 [25]),
    .Y(\soc/cpu/_02037_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06311_  (.A1(\soc/cpu/_02037_ ),
    .A2(\soc/cpu/_02026_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_02038_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_06312_  (.A(\soc/cpu/pcpi_rs2 [26]),
    .B(\soc/cpu/_02038_ ),
    .Y(\soc/cpu/_02039_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_06313_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(\soc/cpu/_02039_ ),
    .Y(\soc/cpu/_02040_ ));
 sky130_fd_sc_hd__a311oi_4 \soc/cpu/_06314_  (.A1(\soc/cpu/_02006_ ),
    .A2(\soc/cpu/_02017_ ),
    .A3(\soc/cpu/_02018_ ),
    .B1(\soc/cpu/_02029_ ),
    .C1(\soc/cpu/_02015_ ),
    .Y(\soc/cpu/_02041_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06315_  (.A(\soc/cpu/_02030_ ),
    .B(\soc/cpu/_02040_ ),
    .C(\soc/cpu/_02041_ ),
    .Y(\soc/cpu/_02042_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06316_  (.A1(\soc/cpu/_02030_ ),
    .A2(\soc/cpu/_02041_ ),
    .B1(\soc/cpu/_02040_ ),
    .Y(\soc/cpu/_02043_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06317_  (.A(net145),
    .B(\soc/cpu/_02043_ ),
    .Y(\soc/cpu/_02044_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06318_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(\soc/cpu/pcpi_rs2 [26]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02045_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06319_  (.A1(\soc/cpu/pcpi_rs1 [26]),
    .A2(\soc/cpu/pcpi_rs2 [26]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_02046_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06320_  (.A1(\soc/cpu/pcpi_rs1 [26]),
    .A2(\soc/cpu/pcpi_rs2 [26]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_02046_ ),
    .Y(\soc/cpu/_02047_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06321_  (.A1(\soc/cpu/_02042_ ),
    .A2(\soc/cpu/_02044_ ),
    .B1(\soc/cpu/_02045_ ),
    .C1(\soc/cpu/_02047_ ),
    .Y(\soc/cpu/alu_out[26] ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06322_  (.A(\soc/cpu/pcpi_rs1 [27]),
    .B(\soc/cpu/pcpi_rs2 [27]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02048_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06323_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(\soc/cpu/pcpi_rs2 [27]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_02049_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06324_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(\soc/cpu/pcpi_rs2 [27]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_02049_ ),
    .Y(\soc/cpu/_02050_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06325_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(\soc/cpu/_02039_ ),
    .Y(\soc/cpu/_02051_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06326_  (.A1(\soc/cpu/_02030_ ),
    .A2(\soc/cpu/_02040_ ),
    .A3(\soc/cpu/_02041_ ),
    .B1(\soc/cpu/_02051_ ),
    .Y(\soc/cpu/_02052_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06327_  (.A(\soc/cpu/pcpi_rs2 [26]),
    .Y(\soc/cpu/_02053_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06328_  (.A(\soc/cpu/_02053_ ),
    .B(\soc/cpu/_02037_ ),
    .C(\soc/cpu/_02026_ ),
    .X(\soc/cpu/_02054_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06329_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_02054_ ),
    .Y(\soc/cpu/_02055_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06330_  (.A(\soc/cpu/pcpi_rs2 [27]),
    .B(\soc/cpu/_02055_ ),
    .Y(\soc/cpu/_02056_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06331_  (.A(\soc/cpu/pcpi_rs1 [27]),
    .B(\soc/cpu/_02056_ ),
    .Y(\soc/cpu/_02057_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_06332_  (.A(\soc/cpu/pcpi_rs1 [27]),
    .B(\soc/cpu/_02056_ ),
    .X(\soc/cpu/_02058_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06333_  (.A(\soc/cpu/_02057_ ),
    .B(\soc/cpu/_02058_ ),
    .X(\soc/cpu/_02059_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06334_  (.A1(\soc/cpu/_02052_ ),
    .A2(\soc/cpu/_02059_ ),
    .B1(\soc/cpu/_01762_ ),
    .Y(\soc/cpu/_02060_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06335_  (.A1(\soc/cpu/_02052_ ),
    .A2(\soc/cpu/_02059_ ),
    .B1(\soc/cpu/_02060_ ),
    .Y(\soc/cpu/_02061_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06336_  (.A(\soc/cpu/_02048_ ),
    .B(\soc/cpu/_02050_ ),
    .C(\soc/cpu/_02061_ ),
    .Y(\soc/cpu/alu_out[27] ));
 sky130_fd_sc_hd__o311ai_4 \soc/cpu/_06337_  (.A1(\soc/cpu/_02030_ ),
    .A2(\soc/cpu/_02040_ ),
    .A3(\soc/cpu/_02041_ ),
    .B1(\soc/cpu/_02057_ ),
    .C1(\soc/cpu/_02051_ ),
    .Y(\soc/cpu/_02062_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06338_  (.A1(\soc/cpu/_01569_ ),
    .A2(\soc/cpu/_02054_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_02063_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06339_  (.A(\soc/cpu/_01568_ ),
    .B(\soc/cpu/_02063_ ),
    .Y(\soc/cpu/_02064_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06340_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .B(\soc/cpu/_02064_ ),
    .X(\soc/cpu/_02065_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06341_  (.A(\soc/cpu/_02065_ ),
    .Y(\soc/cpu/_02066_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06342_  (.A1(\soc/cpu/_02058_ ),
    .A2(\soc/cpu/_02062_ ),
    .B1(\soc/cpu/_02066_ ),
    .Y(\soc/cpu/_02067_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06343_  (.A(\soc/cpu/_02058_ ),
    .B(\soc/cpu/_02066_ ),
    .C(\soc/cpu/_02062_ ),
    .X(\soc/cpu/_02068_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_06344_  (.A(\soc/cpu/_01762_ ),
    .B(\soc/cpu/_02067_ ),
    .C(\soc/cpu/_02068_ ),
    .X(\soc/cpu/_02069_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06345_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .B(\soc/cpu/pcpi_rs2 [28]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02070_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06346_  (.A1(\soc/cpu/pcpi_rs1 [28]),
    .A2(\soc/cpu/pcpi_rs2 [28]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_02071_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06347_  (.A1(\soc/cpu/_01432_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_02069_ ),
    .C1(\soc/cpu/_02070_ ),
    .D1(\soc/cpu/_02071_ ),
    .Y(\soc/cpu/alu_out[28] ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_06348_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .SLEEP(\soc/cpu/_02064_ ),
    .X(\soc/cpu/_02072_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06349_  (.A(\soc/cpu/pcpi_rs2 [28]),
    .B(\soc/cpu/_02063_ ),
    .Y(\soc/cpu/_02073_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06350_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_02073_ ),
    .Y(\soc/cpu/_02074_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06351_  (.A(\soc/cpu/pcpi_rs2 [29]),
    .B(\soc/cpu/_02074_ ),
    .Y(\soc/cpu/_02075_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06352_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(\soc/cpu/_02075_ ),
    .X(\soc/cpu/_02076_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06353_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(\soc/cpu/_02075_ ),
    .Y(\soc/cpu/_02077_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06354_  (.A(\soc/cpu/_02076_ ),
    .B(\soc/cpu/_02077_ ),
    .Y(\soc/cpu/_02078_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06355_  (.A1(\soc/cpu/_02072_ ),
    .A2(\soc/cpu/_02068_ ),
    .B1(\soc/cpu/_02078_ ),
    .Y(\soc/cpu/_02079_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_06356_  (.A(\soc/cpu/_02072_ ),
    .B(\soc/cpu/_02068_ ),
    .C(\soc/cpu/_02078_ ),
    .X(\soc/cpu/_02080_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06357_  (.A(net145),
    .B(\soc/cpu/_02079_ ),
    .C(\soc/cpu/_02080_ ),
    .Y(\soc/cpu/_02081_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06358_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(\soc/cpu/pcpi_rs2 [29]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02082_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06359_  (.A1(\soc/cpu/pcpi_rs1 [29]),
    .A2(\soc/cpu/pcpi_rs2 [29]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_02083_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_06360_  (.A1(\soc/cpu/_01431_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_02081_ ),
    .C1(\soc/cpu/_02082_ ),
    .D1(\soc/cpu/_02083_ ),
    .Y(\soc/cpu/alu_out[29] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06361_  (.A1(\soc/cpu/_01567_ ),
    .A2(\soc/cpu/_02073_ ),
    .B1(\soc/cpu/instr_sub ),
    .Y(\soc/cpu/_02084_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06362_  (.A(\soc/cpu/pcpi_rs2 [30]),
    .B(\soc/cpu/_02084_ ),
    .Y(\soc/cpu/_02085_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06363_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(\soc/cpu/_02085_ ),
    .Y(\soc/cpu/_02086_ ));
 sky130_fd_sc_hd__a311oi_2 \soc/cpu/_06364_  (.A1(\soc/cpu/_02058_ ),
    .A2(\soc/cpu/_02066_ ),
    .A3(\soc/cpu/_02062_ ),
    .B1(\soc/cpu/_02076_ ),
    .C1(\soc/cpu/_02072_ ),
    .Y(\soc/cpu/_02087_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06365_  (.A(\soc/cpu/_02077_ ),
    .B(\soc/cpu/_02086_ ),
    .C(\soc/cpu/_02087_ ),
    .Y(\soc/cpu/_02088_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06366_  (.A1(\soc/cpu/_02077_ ),
    .A2(\soc/cpu/_02087_ ),
    .B1(\soc/cpu/_02086_ ),
    .Y(\soc/cpu/_02089_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06367_  (.A(net145),
    .B(\soc/cpu/_02089_ ),
    .Y(\soc/cpu/_02090_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06368_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(\soc/cpu/pcpi_rs2 [30]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02091_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06369_  (.A1(\soc/cpu/pcpi_rs1 [30]),
    .A2(\soc/cpu/pcpi_rs2 [30]),
    .B1(\soc/cpu/_01759_ ),
    .Y(\soc/cpu/_02092_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06370_  (.A1(\soc/cpu/pcpi_rs1 [30]),
    .A2(\soc/cpu/pcpi_rs2 [30]),
    .B1(\soc/cpu/_01752_ ),
    .B2(\soc/cpu/_02092_ ),
    .Y(\soc/cpu/_02093_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06371_  (.A1(\soc/cpu/_02088_ ),
    .A2(\soc/cpu/_02090_ ),
    .B1(\soc/cpu/_02091_ ),
    .C1(\soc/cpu/_02093_ ),
    .Y(\soc/cpu/alu_out[30] ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_06372_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(\soc/cpu/_02085_ ),
    .X(\soc/cpu/_02094_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06373_  (.A(\soc/cpu/pcpi_rs2 [30]),
    .B(\soc/cpu/_02084_ ),
    .Y(\soc/cpu/_02095_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06374_  (.A(\soc/cpu/instr_sub ),
    .B(\soc/cpu/_02095_ ),
    .Y(\soc/cpu/_02096_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06375_  (.A(\soc/cpu/_01435_ ),
    .B(\soc/cpu/_02096_ ),
    .X(\soc/cpu/_02097_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06376_  (.A1(\soc/cpu/_02094_ ),
    .A2(\soc/cpu/_02088_ ),
    .B1(\soc/cpu/_02097_ ),
    .Y(\soc/cpu/_02098_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_06377_  (.A(\soc/cpu/_02094_ ),
    .B(\soc/cpu/_02088_ ),
    .C(\soc/cpu/_02097_ ),
    .X(\soc/cpu/_02099_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06378_  (.A(\soc/cpu/pcpi_rs1 [31]),
    .B(\soc/cpu/pcpi_rs2 [31]),
    .C(\soc/cpu/_01756_ ),
    .Y(\soc/cpu/_02100_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06379_  (.A1(\soc/cpu/pcpi_rs1 [31]),
    .A2(\soc/cpu/pcpi_rs2 [31]),
    .B1(\soc/cpu/_01752_ ),
    .Y(\soc/cpu/_02101_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06380_  (.A1(\soc/cpu/_01435_ ),
    .A2(\soc/cpu/_01759_ ),
    .B1(\soc/cpu/_02100_ ),
    .C1(\soc/cpu/_02101_ ),
    .Y(\soc/cpu/_02102_ ));
 sky130_fd_sc_hd__a31o_1 \soc/cpu/_06381_  (.A1(net145),
    .A2(\soc/cpu/_02098_ ),
    .A3(\soc/cpu/_02099_ ),
    .B1(\soc/cpu/_02102_ ),
    .X(\soc/cpu/alu_out[31] ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06386_  (.A(\soc/cpu/alu_out_q[0] ),
    .Y(\soc/cpu/_02107_ ));
 sky130_fd_sc_hd__clkinv_4 \soc/cpu/_06387_  (.A(\soc/cpu/latched_branch ),
    .Y(\soc/cpu/_02108_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_06388_  (.A(\soc/cpu/latched_store ),
    .B(\soc/cpu/_02108_ ),
    .Y(\soc/cpu/_02109_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_06390_  (.A1(net297),
    .A2(\soc/cpu/_02107_ ),
    .B1(\soc/cpu/_02109_ ),
    .Y(\soc/cpu/_02111_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06391_  (.A1(net297),
    .A2(net861),
    .B1(\soc/cpu/_02111_ ),
    .Y(\soc/cpu/_02112_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06394_  (.A1(\soc/cpu/reg_next_pc[0] ),
    .A2(\soc/cpu/latched_compr ),
    .B1(\soc/cpu/irq_state[0] ),
    .Y(\soc/cpu/_02115_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_06396_  (.A(\soc/cpu/_00985_ ),
    .B(\soc/cpu/latched_branch ),
    .Y(\soc/cpu/_02117_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_06397_  (.A(\soc/cpu/irq_state[1] ),
    .B(net396),
    .C(\soc/cpu/_02117_ ),
    .Y(\soc/cpu/_02118_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06398_  (.A1(\soc/cpu/irq_state[1] ),
    .A2(\soc/cpu/_00785_ ),
    .B1(\soc/cpu/_02118_ ),
    .B2(\soc/cpu/reg_next_pc[0] ),
    .Y(\soc/cpu/_02119_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_06399_  (.A(\soc/cpu/_02112_ ),
    .B(\soc/cpu/_02115_ ),
    .C(\soc/cpu/_02119_ ),
    .Y(\soc/cpu/cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_06400_  (.A(\soc/cpu/irq_state[1] ),
    .B(\soc/cpu/irq_state[0] ),
    .C(\soc/cpu/_02117_ ),
    .X(\soc/cpu/_02120_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06403_  (.A(net883),
    .B(\soc/cpu/reg_pc[1] ),
    .Y(\soc/cpu/_02123_ ));
 sky130_fd_sc_hd__mux2_2 \soc/cpu/_06404_  (.A0(\soc/cpu/reg_out[1] ),
    .A1(\soc/cpu/alu_out_q[1] ),
    .S(net297),
    .X(\soc/cpu/_02124_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_06405_  (.A1(\soc/cpu/reg_next_pc[1] ),
    .A2(\soc/cpu/irq_state[0] ),
    .B1(\soc/cpu/_02117_ ),
    .B2(\soc/cpu/_02124_ ),
    .C1(\soc/cpu/_00753_ ),
    .C2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02125_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06406_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02123_ ),
    .B1(\soc/cpu/_02125_ ),
    .Y(\soc/cpu/cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__nand2b_2 \soc/cpu/_06408_  (.A_N(\soc/cpu/reg_pc[1] ),
    .B(\soc/cpu/latched_compr ),
    .Y(\soc/cpu/_02127_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06410_  (.A1(\soc/cpu/reg_pc[2] ),
    .A2(\soc/cpu/_02127_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02129_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06411_  (.A1(\soc/cpu/reg_pc[2] ),
    .A2(\soc/cpu/_02127_ ),
    .B1(\soc/cpu/_02129_ ),
    .Y(\soc/cpu/_02130_ ));
 sky130_fd_sc_hd__mux2_4 \soc/cpu/_06413_  (.A0(\soc/cpu/reg_out[2] ),
    .A1(\soc/cpu/alu_out_q[2] ),
    .S(net297),
    .X(\soc/cpu/_02132_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_06414_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[2] ),
    .B1(\soc/cpu/_02117_ ),
    .B2(\soc/cpu/_02132_ ),
    .C1(\soc/cpu/_00762_ ),
    .C2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02133_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_06415_  (.A(\soc/cpu/_02130_ ),
    .B(\soc/cpu/_02133_ ),
    .Y(\soc/cpu/cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06416_  (.A(\soc/cpu/reg_pc[2] ),
    .B(\soc/cpu/_02127_ ),
    .Y(\soc/cpu/_02134_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06417_  (.A(\soc/cpu/reg_pc[3] ),
    .B(\soc/cpu/_02134_ ),
    .X(\soc/cpu/_02135_ ));
 sky130_fd_sc_hd__mux2_2 \soc/cpu/_06418_  (.A0(\soc/cpu/reg_out[3] ),
    .A1(\soc/cpu/alu_out_q[3] ),
    .S(net297),
    .X(\soc/cpu/_02136_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06419_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[3] ),
    .B1(\soc/cpu/_00771_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .X(\soc/cpu/_02137_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06420_  (.A1(\soc/cpu/_02117_ ),
    .A2(\soc/cpu/_02136_ ),
    .B1(\soc/cpu/_02137_ ),
    .Y(\soc/cpu/_02138_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06421_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02135_ ),
    .B1(\soc/cpu/_02138_ ),
    .Y(\soc/cpu/cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_06422_  (.A1(\soc/cpu/reg_pc[2] ),
    .A2(\soc/cpu/reg_pc[3] ),
    .A3(\soc/cpu/_02127_ ),
    .B1(net873),
    .Y(\soc/cpu/_02139_ ));
 sky130_fd_sc_hd__nand4_4 \soc/cpu/_06423_  (.A(\soc/cpu/reg_pc[2] ),
    .B(\soc/cpu/reg_pc[3] ),
    .C(\soc/cpu/reg_pc[4] ),
    .D(\soc/cpu/_02127_ ),
    .Y(\soc/cpu/_02140_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06424_  (.A(\soc/cpu/_02118_ ),
    .B(\soc/cpu/_02140_ ),
    .Y(\soc/cpu/_02141_ ));
 sky130_fd_sc_hd__mux2_2 \soc/cpu/_06425_  (.A0(\soc/cpu/reg_out[4] ),
    .A1(\soc/cpu/alu_out_q[4] ),
    .S(net297),
    .X(\soc/cpu/_02142_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_06426_  (.A(\soc/cpu/irq_state[0] ),
    .Y(\soc/cpu/_02143_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06427_  (.A(\soc/cpu/reg_next_pc[4] ),
    .Y(\soc/cpu/_02144_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06428_  (.A(\soc/cpu/irq_state[1] ),
    .B(\soc/cpu/_00759_ ),
    .Y(\soc/cpu/_02145_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06429_  (.A1(\soc/cpu/_02143_ ),
    .A2(\soc/cpu/_02144_ ),
    .B1(\soc/cpu/_02145_ ),
    .Y(\soc/cpu/_02146_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06430_  (.A1(\soc/cpu/_02117_ ),
    .A2(\soc/cpu/_02142_ ),
    .B1(\soc/cpu/_02146_ ),
    .Y(\soc/cpu/_02147_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06431_  (.A1(\soc/cpu/_02139_ ),
    .A2(\soc/cpu/_02141_ ),
    .B1(\soc/cpu/_02147_ ),
    .Y(\soc/cpu/cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06432_  (.A(\soc/cpu/reg_pc[5] ),
    .B(\soc/cpu/_02140_ ),
    .X(\soc/cpu/_02148_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06436_  (.A0(\soc/cpu/reg_out[5] ),
    .A1(\soc/cpu/alu_out_q[5] ),
    .S(net297),
    .Y(\soc/cpu/_02152_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06437_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02152_ ),
    .Y(\soc/cpu/_02153_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06438_  (.A1(net396),
    .A2(net862),
    .B1(\soc/cpu/_00754_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02153_ ),
    .Y(\soc/cpu/_02154_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06439_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02148_ ),
    .B1(\soc/cpu/_02154_ ),
    .Y(\soc/cpu/cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_06441_  (.A(\soc/cpu/reg_pc[5] ),
    .SLEEP(\soc/cpu/_02140_ ),
    .X(\soc/cpu/_02156_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06442_  (.A1(\soc/cpu/reg_pc[6] ),
    .A2(\soc/cpu/_02156_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02157_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06443_  (.A1(\soc/cpu/reg_pc[6] ),
    .A2(\soc/cpu/_02156_ ),
    .B1(\soc/cpu/_02157_ ),
    .Y(\soc/cpu/_02158_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06444_  (.A0(\soc/cpu/reg_out[6] ),
    .A1(\soc/cpu/alu_out_q[6] ),
    .S(net297),
    .Y(\soc/cpu/_02159_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06445_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02159_ ),
    .Y(\soc/cpu/_02160_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06446_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[6] ),
    .B1(\soc/cpu/_00776_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02160_ ),
    .Y(\soc/cpu/_02161_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_06447_  (.A(\soc/cpu/_02158_ ),
    .B(\soc/cpu/_02161_ ),
    .Y(\soc/cpu/cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06448_  (.A(\soc/cpu/reg_pc[6] ),
    .B(\soc/cpu/_02156_ ),
    .Y(\soc/cpu/_02162_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06449_  (.A(\soc/cpu/reg_pc[7] ),
    .B(\soc/cpu/_02162_ ),
    .X(\soc/cpu/_02163_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06450_  (.A0(\soc/cpu/reg_out[7] ),
    .A1(\soc/cpu/alu_out_q[7] ),
    .S(net297),
    .Y(\soc/cpu/_02164_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06451_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02164_ ),
    .Y(\soc/cpu/_02165_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06452_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[7] ),
    .B1(\soc/cpu/_00758_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02165_ ),
    .Y(\soc/cpu/_02166_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06453_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02163_ ),
    .B1(\soc/cpu/_02166_ ),
    .Y(\soc/cpu/cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_06454_  (.A1(\soc/cpu/reg_pc[6] ),
    .A2(\soc/cpu/reg_pc[7] ),
    .A3(\soc/cpu/_02156_ ),
    .B1(net834),
    .Y(\soc/cpu/_02167_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_06455_  (.A(\soc/cpu/reg_pc[6] ),
    .B(\soc/cpu/reg_pc[7] ),
    .C(\soc/cpu/reg_pc[8] ),
    .D(\soc/cpu/_02156_ ),
    .X(\soc/cpu/_02168_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06457_  (.A0(\soc/cpu/reg_out[8] ),
    .A1(\soc/cpu/alu_out_q[8] ),
    .S(net297),
    .Y(\soc/cpu/_02170_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06458_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02170_ ),
    .Y(\soc/cpu/_02171_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06459_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[8] ),
    .B1(\soc/cpu/_00765_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02171_ ),
    .Y(\soc/cpu/_02172_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_06460_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02167_ ),
    .A3(\soc/cpu/_02168_ ),
    .B1(\soc/cpu/_02172_ ),
    .Y(\soc/cpu/cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06461_  (.A1(\soc/cpu/reg_pc[9] ),
    .A2(\soc/cpu/_02168_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02173_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06462_  (.A1(\soc/cpu/reg_pc[9] ),
    .A2(\soc/cpu/_02168_ ),
    .B1(\soc/cpu/_02173_ ),
    .Y(\soc/cpu/_02174_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06463_  (.A(net396),
    .B(\soc/cpu/reg_next_pc[9] ),
    .Y(\soc/cpu/_02175_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06464_  (.A0(\soc/cpu/reg_out[9] ),
    .A1(\soc/cpu/alu_out_q[9] ),
    .S(net297),
    .X(\soc/cpu/_02176_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06465_  (.A1(\soc/cpu/irq_state[1] ),
    .A2(\soc/cpu/_00774_ ),
    .B1(\soc/cpu/_02117_ ),
    .B2(\soc/cpu/_02176_ ),
    .Y(\soc/cpu/_02177_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_06466_  (.A(\soc/cpu/_02174_ ),
    .B(\soc/cpu/_02175_ ),
    .C(\soc/cpu/_02177_ ),
    .Y(\soc/cpu/cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06467_  (.A(\soc/cpu/reg_pc[9] ),
    .B(\soc/cpu/_02168_ ),
    .Y(\soc/cpu/_02178_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06468_  (.A(\soc/cpu/reg_pc[10] ),
    .B(\soc/cpu/_02178_ ),
    .X(\soc/cpu/_02179_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06469_  (.A0(\soc/cpu/reg_out[10] ),
    .A1(\soc/cpu/alu_out_q[10] ),
    .S(net297),
    .Y(\soc/cpu/_02180_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06470_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02180_ ),
    .Y(\soc/cpu/_02181_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06471_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[10] ),
    .B1(\soc/cpu/_00748_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02181_ ),
    .Y(\soc/cpu/_02182_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06472_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02179_ ),
    .B1(\soc/cpu/_02182_ ),
    .Y(\soc/cpu/cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_06473_  (.A(\soc/cpu/reg_pc[9] ),
    .B(\soc/cpu/reg_pc[10] ),
    .C(\soc/cpu/reg_pc[11] ),
    .D(\soc/cpu/_02168_ ),
    .X(\soc/cpu/_02183_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_06474_  (.A1(\soc/cpu/reg_pc[9] ),
    .A2(\soc/cpu/reg_pc[10] ),
    .A3(\soc/cpu/_02168_ ),
    .B1(\soc/cpu/reg_pc[11] ),
    .Y(\soc/cpu/_02184_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06475_  (.A0(\soc/cpu/reg_out[11] ),
    .A1(\soc/cpu/alu_out_q[11] ),
    .S(net297),
    .Y(\soc/cpu/_02185_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06476_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02185_ ),
    .Y(\soc/cpu/_02186_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06477_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[11] ),
    .B1(\soc/cpu/_00784_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02186_ ),
    .Y(\soc/cpu/_02187_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_06478_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02183_ ),
    .A3(\soc/cpu/_02184_ ),
    .B1(\soc/cpu/_02187_ ),
    .Y(\soc/cpu/cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_06479_  (.A(\soc/cpu/reg_pc[12] ),
    .B(\soc/cpu/_02183_ ),
    .X(\soc/cpu/_02188_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06480_  (.A1(\soc/cpu/reg_pc[12] ),
    .A2(\soc/cpu/_02183_ ),
    .B1(\soc/cpu/_02118_ ),
    .Y(\soc/cpu/_02189_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06481_  (.A0(\soc/cpu/reg_out[12] ),
    .A1(\soc/cpu/alu_out_q[12] ),
    .S(net297),
    .Y(\soc/cpu/_02190_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06482_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02190_ ),
    .Y(\soc/cpu/_02191_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06483_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[12] ),
    .B1(\soc/cpu/_00755_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02191_ ),
    .Y(\soc/cpu/_02192_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06484_  (.A1(\soc/cpu/_02188_ ),
    .A2(\soc/cpu/_02189_ ),
    .B1(\soc/cpu/_02192_ ),
    .Y(\soc/cpu/cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06485_  (.A0(\soc/cpu/reg_out[13] ),
    .A1(\soc/cpu/alu_out_q[13] ),
    .S(net297),
    .Y(\soc/cpu/_02193_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06486_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[13] ),
    .B1(\soc/cpu/_00786_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02194_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06487_  (.A1(\soc/cpu/reg_pc[13] ),
    .A2(\soc/cpu/_02188_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02195_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06488_  (.A1(\soc/cpu/reg_pc[13] ),
    .A2(\soc/cpu/_02188_ ),
    .B1(\soc/cpu/_02195_ ),
    .Y(\soc/cpu/_02196_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_06489_  (.A1(\soc/cpu/_02109_ ),
    .A2(\soc/cpu/_02193_ ),
    .B1(\soc/cpu/_02194_ ),
    .C1(\soc/cpu/_02196_ ),
    .Y(\soc/cpu/cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06490_  (.A1(\soc/cpu/reg_pc[13] ),
    .A2(\soc/cpu/_02188_ ),
    .B1(\soc/cpu/reg_pc[14] ),
    .Y(\soc/cpu/_02197_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06491_  (.A(\soc/cpu/reg_pc[13] ),
    .B(\soc/cpu/reg_pc[14] ),
    .C(\soc/cpu/_02188_ ),
    .X(\soc/cpu/_02198_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_06492_  (.A0(\soc/cpu/reg_out[14] ),
    .A1(\soc/cpu/alu_out_q[14] ),
    .S(net297),
    .Y(\soc/cpu/_02199_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06493_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02199_ ),
    .Y(\soc/cpu/_02200_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06494_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[14] ),
    .B1(\soc/cpu/_00763_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02200_ ),
    .Y(\soc/cpu/_02201_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06495_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02197_ ),
    .A3(\soc/cpu/_02198_ ),
    .B1(\soc/cpu/_02201_ ),
    .Y(\soc/cpu/cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_06496_  (.A(\soc/cpu/reg_pc[15] ),
    .B(\soc/cpu/_02198_ ),
    .X(\soc/cpu/_02202_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06497_  (.A1(\soc/cpu/reg_pc[15] ),
    .A2(\soc/cpu/_02198_ ),
    .B1(\soc/cpu/_02118_ ),
    .Y(\soc/cpu/_02203_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06498_  (.A0(\soc/cpu/reg_out[15] ),
    .A1(\soc/cpu/alu_out_q[15] ),
    .S(net297),
    .Y(\soc/cpu/_02204_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06499_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02204_ ),
    .Y(\soc/cpu/_02205_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06500_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[15] ),
    .B1(\soc/cpu/_00773_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02205_ ),
    .Y(\soc/cpu/_02206_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06501_  (.A1(\soc/cpu/_02202_ ),
    .A2(\soc/cpu/_02203_ ),
    .B1(\soc/cpu/_02206_ ),
    .Y(\soc/cpu/cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06502_  (.A0(\soc/cpu/reg_out[16] ),
    .A1(\soc/cpu/alu_out_q[16] ),
    .S(net297),
    .Y(\soc/cpu/_02207_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06503_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[16] ),
    .B1(\soc/cpu/_00781_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02208_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06504_  (.A1(\soc/cpu/reg_pc[16] ),
    .A2(\soc/cpu/_02202_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02209_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06505_  (.A1(\soc/cpu/reg_pc[16] ),
    .A2(\soc/cpu/_02202_ ),
    .B1(\soc/cpu/_02209_ ),
    .Y(\soc/cpu/_02210_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_06506_  (.A1(\soc/cpu/_02109_ ),
    .A2(\soc/cpu/_02207_ ),
    .B1(\soc/cpu/_02208_ ),
    .C1(\soc/cpu/_02210_ ),
    .Y(\soc/cpu/cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_06507_  (.A(\soc/cpu/reg_pc[16] ),
    .B(\soc/cpu/reg_pc[17] ),
    .C(\soc/cpu/_02202_ ),
    .X(\soc/cpu/_02211_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06508_  (.A1(\soc/cpu/reg_pc[16] ),
    .A2(\soc/cpu/_02202_ ),
    .B1(\soc/cpu/reg_pc[17] ),
    .Y(\soc/cpu/_02212_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06509_  (.A0(\soc/cpu/reg_out[17] ),
    .A1(\soc/cpu/alu_out_q[17] ),
    .S(net297),
    .Y(\soc/cpu/_02213_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06510_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02213_ ),
    .Y(\soc/cpu/_02214_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06511_  (.A1(net396),
    .A2(\soc/cpu/reg_next_pc[17] ),
    .B1(\soc/cpu/_00770_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02214_ ),
    .Y(\soc/cpu/_02215_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_06512_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02211_ ),
    .A3(\soc/cpu/_02212_ ),
    .B1(\soc/cpu/_02215_ ),
    .Y(\soc/cpu/cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_06513_  (.A(\soc/cpu/reg_pc[18] ),
    .B(\soc/cpu/_02211_ ),
    .X(\soc/cpu/_02216_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06514_  (.A1(\soc/cpu/reg_pc[18] ),
    .A2(\soc/cpu/_02211_ ),
    .B1(\soc/cpu/_02118_ ),
    .Y(\soc/cpu/_02217_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06515_  (.A0(\soc/cpu/reg_out[18] ),
    .A1(\soc/cpu/alu_out_q[18] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02218_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06516_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02218_ ),
    .Y(\soc/cpu/_02219_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06517_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[18] ),
    .B1(\soc/cpu/_00750_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02219_ ),
    .Y(\soc/cpu/_02220_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06518_  (.A1(\soc/cpu/_02216_ ),
    .A2(\soc/cpu/_02217_ ),
    .B1(\soc/cpu/_02220_ ),
    .Y(\soc/cpu/cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06519_  (.A1(\soc/cpu/reg_pc[19] ),
    .A2(\soc/cpu/_02216_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02221_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06520_  (.A1(\soc/cpu/reg_pc[19] ),
    .A2(\soc/cpu/_02216_ ),
    .B1(\soc/cpu/_02221_ ),
    .Y(\soc/cpu/_02222_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06521_  (.A0(\soc/cpu/reg_out[19] ),
    .A1(\soc/cpu/alu_out_q[19] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02223_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06522_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02223_ ),
    .Y(\soc/cpu/_02224_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06523_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[19] ),
    .B1(\soc/cpu/_00779_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02224_ ),
    .Y(\soc/cpu/_02225_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_06524_  (.A(\soc/cpu/_02222_ ),
    .B(\soc/cpu/_02225_ ),
    .Y(\soc/cpu/cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06525_  (.A1(\soc/cpu/reg_pc[19] ),
    .A2(\soc/cpu/_02216_ ),
    .B1(\soc/cpu/reg_pc[20] ),
    .Y(\soc/cpu/_02226_ ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_06526_  (.A(\soc/cpu/reg_pc[19] ),
    .B(\soc/cpu/reg_pc[20] ),
    .C(\soc/cpu/_02216_ ),
    .X(\soc/cpu/_02227_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06527_  (.A0(\soc/cpu/reg_out[20] ),
    .A1(\soc/cpu/alu_out_q[20] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02228_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06528_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02228_ ),
    .Y(\soc/cpu/_02229_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06529_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[20] ),
    .B1(\soc/cpu/_00749_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02229_ ),
    .Y(\soc/cpu/_02230_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_06530_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02226_ ),
    .A3(\soc/cpu/_02227_ ),
    .B1(\soc/cpu/_02230_ ),
    .Y(\soc/cpu/cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06531_  (.A0(\soc/cpu/reg_out[21] ),
    .A1(\soc/cpu/alu_out_q[21] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02231_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06532_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[21] ),
    .B1(\soc/cpu/_00764_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02232_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06533_  (.A1(\soc/cpu/reg_pc[21] ),
    .A2(\soc/cpu/_02227_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02233_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06534_  (.A1(\soc/cpu/reg_pc[21] ),
    .A2(\soc/cpu/_02227_ ),
    .B1(\soc/cpu/_02233_ ),
    .Y(\soc/cpu/_02234_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_06535_  (.A1(\soc/cpu/_02109_ ),
    .A2(\soc/cpu/_02231_ ),
    .B1(\soc/cpu/_02232_ ),
    .C1(\soc/cpu/_02234_ ),
    .Y(\soc/cpu/cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06536_  (.A1(\soc/cpu/reg_pc[21] ),
    .A2(\soc/cpu/_02227_ ),
    .B1(\soc/cpu/reg_pc[22] ),
    .Y(\soc/cpu/_02235_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06537_  (.A(\soc/cpu/reg_pc[21] ),
    .B(\soc/cpu/reg_pc[22] ),
    .C(\soc/cpu/_02227_ ),
    .X(\soc/cpu/_02236_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06538_  (.A0(\soc/cpu/reg_out[22] ),
    .A1(\soc/cpu/alu_out_q[22] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02237_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06539_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02237_ ),
    .Y(\soc/cpu/_02238_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_06540_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[22] ),
    .B1(\soc/cpu/_00783_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02238_ ),
    .Y(\soc/cpu/_02239_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06541_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02235_ ),
    .A3(\soc/cpu/_02236_ ),
    .B1(\soc/cpu/_02239_ ),
    .Y(\soc/cpu/cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_06542_  (.A(\soc/cpu/reg_pc[23] ),
    .B(\soc/cpu/_02236_ ),
    .X(\soc/cpu/_02240_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06543_  (.A1(\soc/cpu/reg_pc[23] ),
    .A2(\soc/cpu/_02236_ ),
    .B1(\soc/cpu/_02118_ ),
    .Y(\soc/cpu/_02241_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06544_  (.A0(\soc/cpu/reg_out[23] ),
    .A1(\soc/cpu/alu_out_q[23] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02242_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06545_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02242_ ),
    .Y(\soc/cpu/_02243_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06546_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[23] ),
    .B1(\soc/cpu/_00768_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02243_ ),
    .Y(\soc/cpu/_02244_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06547_  (.A1(\soc/cpu/_02240_ ),
    .A2(\soc/cpu/_02241_ ),
    .B1(\soc/cpu/_02244_ ),
    .Y(\soc/cpu/cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06548_  (.A0(\soc/cpu/reg_out[24] ),
    .A1(\soc/cpu/alu_out_q[24] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02245_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06549_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[24] ),
    .B1(\soc/cpu/_00780_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02246_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06550_  (.A1(\soc/cpu/reg_pc[24] ),
    .A2(\soc/cpu/_02240_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02247_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06551_  (.A1(\soc/cpu/reg_pc[24] ),
    .A2(\soc/cpu/_02240_ ),
    .B1(\soc/cpu/_02247_ ),
    .Y(\soc/cpu/_02248_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_06552_  (.A1(\soc/cpu/_02109_ ),
    .A2(\soc/cpu/_02245_ ),
    .B1(\soc/cpu/_02246_ ),
    .C1(\soc/cpu/_02248_ ),
    .Y(\soc/cpu/cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06553_  (.A1(\soc/cpu/reg_pc[24] ),
    .A2(\soc/cpu/_02240_ ),
    .B1(\soc/cpu/reg_pc[25] ),
    .Y(\soc/cpu/_02249_ ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_06554_  (.A(\soc/cpu/reg_pc[24] ),
    .B(\soc/cpu/reg_pc[25] ),
    .C(\soc/cpu/_02240_ ),
    .X(\soc/cpu/_02250_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_06555_  (.A0(\soc/cpu/reg_out[25] ),
    .A1(\soc/cpu/alu_out_q[25] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02251_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06556_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02251_ ),
    .Y(\soc/cpu/_02252_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06557_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[25] ),
    .B1(\soc/cpu/_00752_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02252_ ),
    .Y(\soc/cpu/_02253_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_06558_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02249_ ),
    .A3(\soc/cpu/_02250_ ),
    .B1(\soc/cpu/_02253_ ),
    .Y(\soc/cpu/cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06559_  (.A0(\soc/cpu/reg_out[26] ),
    .A1(\soc/cpu/alu_out_q[26] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02254_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06560_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[26] ),
    .B1(\soc/cpu/_00775_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02255_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06561_  (.A1(\soc/cpu/reg_pc[26] ),
    .A2(\soc/cpu/_02250_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02256_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06562_  (.A1(\soc/cpu/reg_pc[26] ),
    .A2(\soc/cpu/_02250_ ),
    .B1(\soc/cpu/_02256_ ),
    .Y(\soc/cpu/_02257_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_06563_  (.A1(\soc/cpu/_02109_ ),
    .A2(\soc/cpu/_02254_ ),
    .B1(\soc/cpu/_02255_ ),
    .C1(\soc/cpu/_02257_ ),
    .Y(\soc/cpu/cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_06564_  (.A(\soc/cpu/reg_pc[26] ),
    .B(\soc/cpu/reg_pc[27] ),
    .C(\soc/cpu/_02250_ ),
    .X(\soc/cpu/_02258_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06565_  (.A1(\soc/cpu/reg_pc[26] ),
    .A2(\soc/cpu/_02250_ ),
    .B1(\soc/cpu/reg_pc[27] ),
    .Y(\soc/cpu/_02259_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_06566_  (.A0(\soc/cpu/reg_out[27] ),
    .A1(\soc/cpu/alu_out_q[27] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02260_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06567_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02260_ ),
    .Y(\soc/cpu/_02261_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_06568_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[27] ),
    .B1(\soc/cpu/_00760_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02261_ ),
    .Y(\soc/cpu/_02262_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06569_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02258_ ),
    .A3(\soc/cpu/_02259_ ),
    .B1(\soc/cpu/_02262_ ),
    .Y(\soc/cpu/cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_06570_  (.A0(\soc/cpu/reg_out[28] ),
    .A1(\soc/cpu/alu_out_q[28] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02263_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06571_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[28] ),
    .B1(\soc/cpu/_00757_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_02264_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06572_  (.A1(\soc/cpu/reg_pc[28] ),
    .A2(\soc/cpu/_02258_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02265_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06573_  (.A1(\soc/cpu/reg_pc[28] ),
    .A2(\soc/cpu/_02258_ ),
    .B1(\soc/cpu/_02265_ ),
    .Y(\soc/cpu/_02266_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_06574_  (.A1(\soc/cpu/_02109_ ),
    .A2(\soc/cpu/_02263_ ),
    .B1(\soc/cpu/_02264_ ),
    .C1(\soc/cpu/_02266_ ),
    .Y(\soc/cpu/cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_06575_  (.A(\soc/cpu/reg_pc[28] ),
    .B(\soc/cpu/reg_pc[29] ),
    .C(\soc/cpu/_02258_ ),
    .X(\soc/cpu/_02267_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06576_  (.A1(\soc/cpu/reg_pc[28] ),
    .A2(\soc/cpu/_02258_ ),
    .B1(\soc/cpu/reg_pc[29] ),
    .Y(\soc/cpu/_02268_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_06577_  (.A0(\soc/cpu/reg_out[29] ),
    .A1(\soc/cpu/alu_out_q[29] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02269_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06578_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02269_ ),
    .Y(\soc/cpu/_02270_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06579_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[29] ),
    .B1(\soc/cpu/_00747_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02270_ ),
    .Y(\soc/cpu/_02271_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_06580_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02267_ ),
    .A3(\soc/cpu/_02268_ ),
    .B1(\soc/cpu/_02271_ ),
    .Y(\soc/cpu/cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06581_  (.A1(\soc/cpu/reg_pc[30] ),
    .A2(\soc/cpu/_02267_ ),
    .B1(\soc/cpu/_02120_ ),
    .Y(\soc/cpu/_02272_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06582_  (.A1(\soc/cpu/reg_pc[30] ),
    .A2(\soc/cpu/_02267_ ),
    .B1(\soc/cpu/_02272_ ),
    .Y(\soc/cpu/_02273_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_06583_  (.A0(\soc/cpu/reg_out[30] ),
    .A1(\soc/cpu/alu_out_q[30] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02274_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06584_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02274_ ),
    .Y(\soc/cpu/_02275_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06585_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[30] ),
    .B1(\soc/cpu/_00769_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02275_ ),
    .Y(\soc/cpu/_02276_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_06586_  (.A(\soc/cpu/_02273_ ),
    .B(\soc/cpu/_02276_ ),
    .Y(\soc/cpu/cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06587_  (.A(\soc/cpu/reg_pc[30] ),
    .B(\soc/cpu/_02267_ ),
    .Y(\soc/cpu/_02277_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_06588_  (.A(\soc/cpu/reg_pc[31] ),
    .B(\soc/cpu/_02277_ ),
    .X(\soc/cpu/_02278_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_06589_  (.A0(\soc/cpu/reg_out[31] ),
    .A1(\soc/cpu/alu_out_q[31] ),
    .S(\soc/cpu/latched_stalu ),
    .Y(\soc/cpu/_02279_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06590_  (.A(\soc/cpu/_02109_ ),
    .B(\soc/cpu/_02279_ ),
    .Y(\soc/cpu/_02280_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06591_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/reg_next_pc[31] ),
    .B1(\soc/cpu/_00778_ ),
    .B2(\soc/cpu/irq_state[1] ),
    .C1(\soc/cpu/_02280_ ),
    .Y(\soc/cpu/_02281_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06592_  (.A1(\soc/cpu/_02120_ ),
    .A2(\soc/cpu/_02278_ ),
    .B1(\soc/cpu/_02281_ ),
    .Y(\soc/cpu/cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06593_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02282_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06594_  (.A_N(\soc/cpu/mem_wordsize[2] ),
    .B(\soc/cpu/mem_wordsize[1] ),
    .Y(\soc/cpu/_02283_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06595_  (.A(\soc/cpu/_02282_ ),
    .B(\soc/cpu/_02283_ ),
    .Y(\soc/cpu/_02284_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_06596_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/pcpi_rs1 [1]),
    .B1(\soc/cpu/_02284_ ),
    .Y(\soc/cpu/mem_la_wstrb [0]));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06597_  (.A1(\soc/cpu/_01490_ ),
    .A2(\soc/cpu/pcpi_rs1 [1]),
    .B1(\soc/cpu/_02284_ ),
    .Y(\soc/cpu/mem_la_wstrb [1]));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_06598_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .SLEEP(\soc/cpu/pcpi_rs1 [0]),
    .X(\soc/cpu/_02285_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06599_  (.A1(\soc/cpu/mem_wordsize[2] ),
    .A2(\soc/cpu/mem_wordsize[1] ),
    .B1(\soc/cpu/_02282_ ),
    .Y(\soc/cpu/_02286_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_06600_  (.A(\soc/cpu/_02285_ ),
    .B(\soc/cpu/_02286_ ),
    .X(\soc/cpu/mem_la_wstrb [2]));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_06601_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/pcpi_rs1 [1]),
    .B1(\soc/cpu/_02286_ ),
    .X(\soc/cpu/mem_la_wstrb [3]));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06602_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/mem_la_wdata [0]),
    .B1(net780),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02287_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06603_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01845_ ),
    .B1(\soc/cpu/_02287_ ),
    .Y(\soc/cpu/mem_la_wdata [8]));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06604_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/mem_la_wdata [1]),
    .B1(net781),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02288_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06605_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01538_ ),
    .B1(\soc/cpu/_02288_ ),
    .Y(\soc/cpu/mem_la_wdata [9]));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06606_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/mem_la_wdata [2]),
    .B1(\soc/cpu/pcpi_rs2 [10]),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02289_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06607_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01869_ ),
    .B1(\soc/cpu/_02289_ ),
    .Y(\soc/cpu/mem_la_wdata [10]));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06608_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/mem_la_wdata [3]),
    .B1(net777),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02290_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06609_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01537_ ),
    .B1(\soc/cpu/_02290_ ),
    .Y(\soc/cpu/mem_la_wdata [11]));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06610_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/mem_la_wdata [4]),
    .B1(\soc/cpu/pcpi_rs2 [12]),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02291_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06611_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01534_ ),
    .B1(\soc/cpu/_02291_ ),
    .Y(\soc/cpu/mem_la_wdata [12]));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06612_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/mem_la_wdata [5]),
    .B1(\soc/cpu/pcpi_rs2 [13]),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02292_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06613_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01533_ ),
    .B1(\soc/cpu/_02292_ ),
    .Y(\soc/cpu/mem_la_wdata [13]));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_06614_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(net776),
    .B1(\soc/cpu/pcpi_rs2 [14]),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_02293_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_06615_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01912_ ),
    .B1(\soc/cpu/_02293_ ),
    .Y(\soc/cpu/mem_la_wdata [14]));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06616_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(net773),
    .B1(\soc/cpu/pcpi_rs2 [15]),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .X(\soc/cpu/_02294_ ));
 sky130_fd_sc_hd__o21bai_2 \soc/cpu/_06617_  (.A1(\soc/cpu/mem_wordsize[1] ),
    .A2(\soc/cpu/_01530_ ),
    .B1_N(\soc/cpu/_02294_ ),
    .Y(\soc/cpu/mem_la_wdata [15]));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_06618_  (.A(\soc/cpu/mem_wordsize[2] ),
    .B(\soc/cpu/mem_wordsize[1] ),
    .Y(\soc/cpu/_02295_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06619_  (.A0(\soc/cpu/mem_la_wdata [0]),
    .A1(\soc/cpu/pcpi_rs2 [16]),
    .S(net157),
    .X(\soc/cpu/mem_la_wdata [16]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06622_  (.A(\soc/cpu/pcpi_rs2 [17]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02298_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06623_  (.A1(\soc/cpu/_01521_ ),
    .A2(net157),
    .B1(\soc/cpu/_02298_ ),
    .Y(\soc/cpu/mem_la_wdata [17]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06624_  (.A(\soc/cpu/pcpi_rs2 [18]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02299_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06625_  (.A1(\soc/cpu/_01520_ ),
    .A2(net157),
    .B1(\soc/cpu/_02299_ ),
    .Y(\soc/cpu/mem_la_wdata [18]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06626_  (.A(\soc/cpu/pcpi_rs2 [19]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02300_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06627_  (.A1(\soc/cpu/_01519_ ),
    .A2(net157),
    .B1(\soc/cpu/_02300_ ),
    .Y(\soc/cpu/mem_la_wdata [19]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06628_  (.A(\soc/cpu/pcpi_rs2 [20]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02301_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06629_  (.A1(\soc/cpu/_01518_ ),
    .A2(net157),
    .B1(\soc/cpu/_02301_ ),
    .Y(\soc/cpu/mem_la_wdata [20]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06630_  (.A(\soc/cpu/pcpi_rs2 [21]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02302_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06631_  (.A1(\soc/cpu/_01517_ ),
    .A2(net157),
    .B1(\soc/cpu/_02302_ ),
    .Y(\soc/cpu/mem_la_wdata [21]));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06632_  (.A0(net776),
    .A1(net754),
    .S(\soc/cpu/_02295_ ),
    .X(\soc/cpu/mem_la_wdata [22]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06634_  (.A(\soc/cpu/pcpi_rs2 [23]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02304_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_06635_  (.A1(\soc/cpu/_01516_ ),
    .A2(\soc/cpu/_02295_ ),
    .B1(\soc/cpu/_02304_ ),
    .Y(\soc/cpu/mem_la_wdata [23]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06637_  (.A(\soc/cpu/pcpi_rs2 [24]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02306_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06638_  (.A(\soc/cpu/_02287_ ),
    .B(\soc/cpu/_02306_ ),
    .Y(\soc/cpu/mem_la_wdata [24]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06639_  (.A(\soc/cpu/pcpi_rs2 [25]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02307_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06640_  (.A(\soc/cpu/_02288_ ),
    .B(\soc/cpu/_02307_ ),
    .Y(\soc/cpu/mem_la_wdata [25]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06641_  (.A(\soc/cpu/pcpi_rs2 [26]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02308_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06642_  (.A(\soc/cpu/_02289_ ),
    .B(\soc/cpu/_02308_ ),
    .Y(\soc/cpu/mem_la_wdata [26]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06643_  (.A(\soc/cpu/pcpi_rs2 [27]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02309_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06644_  (.A(\soc/cpu/_02290_ ),
    .B(\soc/cpu/_02309_ ),
    .Y(\soc/cpu/mem_la_wdata [27]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06645_  (.A(\soc/cpu/pcpi_rs2 [28]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02310_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06646_  (.A(\soc/cpu/_02291_ ),
    .B(\soc/cpu/_02310_ ),
    .Y(\soc/cpu/mem_la_wdata [28]));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_06647_  (.A(\soc/cpu/pcpi_rs2 [29]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02311_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06648_  (.A(\soc/cpu/_02292_ ),
    .B(\soc/cpu/_02311_ ),
    .Y(\soc/cpu/mem_la_wdata [29]));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06649_  (.A(\soc/cpu/pcpi_rs2 [30]),
    .B(\soc/cpu/_02295_ ),
    .Y(\soc/cpu/_02312_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06650_  (.A(\soc/cpu/_02293_ ),
    .B(\soc/cpu/_02312_ ),
    .Y(\soc/cpu/mem_la_wdata [30]));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_06651_  (.A1(\soc/cpu/pcpi_rs2 [31]),
    .A2(\soc/cpu/_02295_ ),
    .B1(\soc/cpu/_02294_ ),
    .X(\soc/cpu/mem_la_wdata [31]));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/_06652_  (.A1(\soc/cpu/irq_pending[1] ),
    .A2(\soc/cpu/_00935_ ),
    .B1(\soc/cpu/_00992_ ),
    .B2(\soc/cpu/irq_mask[1] ),
    .C1(_074_),
    .Y(\soc/cpu/_02313_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06653_  (.A_N(net419),
    .B(\soc/cpu/_02313_ ),
    .Y(\soc/cpu/_00012_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06656_  (.A1(\soc/cpu/irq_mask[3] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[3] ),
    .Y(\soc/cpu/_02316_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06657_  (.A1(net132),
    .A2(\soc/cpu/_02316_ ),
    .B1_N(net420),
    .Y(\soc/cpu/_00026_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06658_  (.A1(\soc/cpu/irq_mask[4] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[4] ),
    .Y(\soc/cpu/_02317_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06659_  (.A1(net131),
    .A2(\soc/cpu/_02317_ ),
    .B1_N(net421),
    .Y(\soc/cpu/_00027_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06661_  (.A1(\soc/cpu/irq_mask[5] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[5] ),
    .Y(\soc/cpu/_02319_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06662_  (.A1(net132),
    .A2(\soc/cpu/_02319_ ),
    .B1_N(net416),
    .Y(\soc/cpu/_00028_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06663_  (.A1(\soc/cpu/irq_mask[6] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[6] ),
    .Y(\soc/cpu/_02320_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06664_  (.A1(net132),
    .A2(\soc/cpu/_02320_ ),
    .B1_N(net417),
    .Y(\soc/cpu/_00029_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06665_  (.A1(\soc/cpu/irq_mask[7] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[7] ),
    .Y(\soc/cpu/_02321_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06666_  (.A1(net132),
    .A2(\soc/cpu/_02321_ ),
    .B1_N(net418),
    .Y(\soc/cpu/_00030_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06667_  (.A1(\soc/cpu/irq_mask[8] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[8] ),
    .Y(\soc/cpu/_02322_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06668_  (.A1(net131),
    .A2(\soc/cpu/_02322_ ),
    .B1_N(net422),
    .Y(\soc/cpu/_00031_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06669_  (.A1(\soc/cpu/irq_mask[9] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[9] ),
    .Y(\soc/cpu/_02323_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06670_  (.A1(net131),
    .A2(\soc/cpu/_02323_ ),
    .B1_N(net423),
    .Y(\soc/cpu/_00032_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06671_  (.A1(\soc/cpu/irq_mask[10] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[10] ),
    .Y(\soc/cpu/_02324_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06672_  (.A1(net131),
    .A2(\soc/cpu/_02324_ ),
    .B1_N(net424),
    .Y(\soc/cpu/_00002_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06674_  (.A1(net887),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[11] ),
    .Y(\soc/cpu/_02326_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06675_  (.A1(net131),
    .A2(\soc/cpu/_02326_ ),
    .B1_N(net425),
    .Y(\soc/cpu/_00003_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06676_  (.A1(\soc/cpu/irq_mask[12] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[12] ),
    .Y(\soc/cpu/_02327_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06677_  (.A1(net131),
    .A2(\soc/cpu/_02327_ ),
    .B1_N(net426),
    .Y(\soc/cpu/_00004_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06678_  (.A1(\soc/cpu/irq_mask[13] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[13] ),
    .Y(\soc/cpu/_02328_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06679_  (.A1(net131),
    .A2(\soc/cpu/_02328_ ),
    .B1_N(net427),
    .Y(\soc/cpu/_00005_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06680_  (.A1(\soc/cpu/irq_mask[14] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[14] ),
    .Y(\soc/cpu/_02329_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06681_  (.A1(net131),
    .A2(\soc/cpu/_02329_ ),
    .B1_N(net428),
    .Y(\soc/cpu/_00006_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06683_  (.A1(\soc/cpu/irq_mask[15] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[15] ),
    .Y(\soc/cpu/_02331_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06684_  (.A1(net131),
    .A2(\soc/cpu/_02331_ ),
    .B1_N(net429),
    .Y(\soc/cpu/_00007_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06685_  (.A1(\soc/cpu/irq_mask[16] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[16] ),
    .Y(\soc/cpu/_02332_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06686_  (.A1(net131),
    .A2(\soc/cpu/_02332_ ),
    .B1_N(net430),
    .Y(\soc/cpu/_00008_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06687_  (.A1(\soc/cpu/irq_mask[17] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[17] ),
    .Y(\soc/cpu/_02333_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06688_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02333_ ),
    .B1_N(net431),
    .Y(\soc/cpu/_00009_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06689_  (.A1(net866),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[18] ),
    .Y(\soc/cpu/_02334_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06690_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02334_ ),
    .B1_N(net432),
    .Y(\soc/cpu/_00010_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06691_  (.A1(\soc/cpu/irq_mask[19] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[19] ),
    .Y(\soc/cpu/_02335_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06692_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02335_ ),
    .B1_N(net433),
    .Y(\soc/cpu/_00011_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06693_  (.A1(\soc/cpu/irq_mask[20] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[20] ),
    .Y(\soc/cpu/_02336_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06694_  (.A1(net131),
    .A2(\soc/cpu/_02336_ ),
    .B1_N(net434),
    .Y(\soc/cpu/_00013_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06696_  (.A1(\soc/cpu/irq_mask[21] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[21] ),
    .Y(\soc/cpu/_02338_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06697_  (.A1(net131),
    .A2(\soc/cpu/_02338_ ),
    .B1_N(net435),
    .Y(\soc/cpu/_00014_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06698_  (.A1(\soc/cpu/irq_mask[22] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[22] ),
    .Y(\soc/cpu/_02339_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06699_  (.A1(net131),
    .A2(\soc/cpu/_02339_ ),
    .B1_N(net436),
    .Y(\soc/cpu/_00015_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06700_  (.A1(\soc/cpu/irq_mask[23] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[23] ),
    .Y(\soc/cpu/_02340_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06701_  (.A1(net131),
    .A2(\soc/cpu/_02340_ ),
    .B1_N(net437),
    .Y(\soc/cpu/_00016_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06702_  (.A1(\soc/cpu/irq_mask[24] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[24] ),
    .Y(\soc/cpu/_02341_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06703_  (.A1(net131),
    .A2(\soc/cpu/_02341_ ),
    .B1_N(net438),
    .Y(\soc/cpu/_00017_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06705_  (.A1(\soc/cpu/irq_mask[25] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[25] ),
    .Y(\soc/cpu/_02343_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06706_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02343_ ),
    .B1_N(net439),
    .Y(\soc/cpu/_00018_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06707_  (.A1(\soc/cpu/irq_mask[26] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[26] ),
    .Y(\soc/cpu/_02344_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06708_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02344_ ),
    .B1_N(net440),
    .Y(\soc/cpu/_00019_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06709_  (.A1(\soc/cpu/irq_mask[27] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[27] ),
    .Y(\soc/cpu/_02345_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06710_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02345_ ),
    .B1_N(net441),
    .Y(\soc/cpu/_00020_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06711_  (.A1(\soc/cpu/irq_mask[28] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[28] ),
    .Y(\soc/cpu/_02346_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06712_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02346_ ),
    .B1_N(net442),
    .Y(\soc/cpu/_00021_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06713_  (.A1(\soc/cpu/irq_mask[29] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[29] ),
    .Y(\soc/cpu/_02347_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06714_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02347_ ),
    .B1_N(net443),
    .Y(\soc/cpu/_00022_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06715_  (.A1(\soc/cpu/irq_mask[30] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[30] ),
    .Y(\soc/cpu/_02348_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06716_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02348_ ),
    .B1_N(net444),
    .Y(\soc/cpu/_00024_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06717_  (.A1(\soc/cpu/irq_mask[31] ),
    .A2(\soc/cpu/_00992_ ),
    .B1(\soc/cpu/irq_pending[31] ),
    .Y(\soc/cpu/_02349_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_06718_  (.A1(\soc/cpu/_00840_ ),
    .A2(\soc/cpu/_02349_ ),
    .B1_N(net445),
    .Y(\soc/cpu/_00025_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06719_  (.A_N(\soc/cpu/mem_state[1] ),
    .B(net892),
    .Y(\soc/cpu/_02350_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06720_  (.A(\soc/cpu/_00721_ ),
    .B(\soc/cpu/_02350_ ),
    .Y(\soc/cpu/_02351_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_06721_  (.A(net132),
    .B(\soc/cpu/trap ),
    .Y(\soc/cpu/_02352_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06722_  (.A(\soc/mem_rdata[0] ),
    .B(\soc/mem_rdata[1] ),
    .Y(\soc/cpu/_02353_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06723_  (.A(\soc/cpu/mem_do_rdata ),
    .B(\soc/cpu/mem_la_read ),
    .Y(\soc/cpu/_02354_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06724_  (.A1(\soc/cpu/mem_la_secondword ),
    .A2(\soc/cpu/_02353_ ),
    .B1(\soc/cpu/_02354_ ),
    .Y(\soc/cpu/_02355_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06725_  (.A1(\soc/cpu/_00715_ ),
    .A2(\soc/cpu/_00745_ ),
    .B1(\soc/cpu/_02355_ ),
    .Y(\soc/cpu/_02356_ ));
 sky130_fd_sc_hd__and3_4 \soc/cpu/_06726_  (.A(\soc/cpu/_02351_ ),
    .B(\soc/cpu/_02352_ ),
    .C(\soc/cpu/_02356_ ),
    .X(\soc/cpu/_02357_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06729_  (.A0(\soc/cpu/mem_16bit_buffer[0] ),
    .A1(\soc/mem_rdata[16] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00082_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06730_  (.A0(\soc/cpu/mem_16bit_buffer[1] ),
    .A1(\soc/mem_rdata[17] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00083_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06731_  (.A0(\soc/cpu/mem_16bit_buffer[2] ),
    .A1(\soc/mem_rdata[18] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00084_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06732_  (.A0(\soc/cpu/mem_16bit_buffer[3] ),
    .A1(\soc/mem_rdata[19] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00085_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06733_  (.A0(\soc/cpu/mem_16bit_buffer[4] ),
    .A1(\soc/mem_rdata[20] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00086_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06734_  (.A0(\soc/cpu/mem_16bit_buffer[5] ),
    .A1(\soc/mem_rdata[21] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00087_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06735_  (.A0(\soc/cpu/mem_16bit_buffer[6] ),
    .A1(\soc/mem_rdata[22] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00088_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06736_  (.A0(\soc/cpu/mem_16bit_buffer[7] ),
    .A1(\soc/mem_rdata[23] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00089_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06737_  (.A0(\soc/cpu/mem_16bit_buffer[8] ),
    .A1(\soc/mem_rdata[24] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00090_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06738_  (.A0(\soc/cpu/mem_16bit_buffer[9] ),
    .A1(\soc/mem_rdata[25] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00091_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06739_  (.A0(\soc/cpu/mem_16bit_buffer[10] ),
    .A1(\soc/mem_rdata[26] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00092_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06740_  (.A0(\soc/cpu/mem_16bit_buffer[11] ),
    .A1(\soc/mem_rdata[27] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00093_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06741_  (.A0(\soc/cpu/mem_16bit_buffer[12] ),
    .A1(\soc/mem_rdata[28] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00094_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06742_  (.A0(\soc/cpu/mem_16bit_buffer[13] ),
    .A1(\soc/mem_rdata[29] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00095_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06743_  (.A0(\soc/cpu/mem_16bit_buffer[14] ),
    .A1(\soc/mem_rdata[30] ),
    .S(\soc/cpu/_02357_ ),
    .X(\soc/cpu/_00096_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06744_  (.A(\soc/mem_rdata[31] ),
    .Y(\soc/cpu/_02360_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06745_  (.A(\soc/cpu/mem_16bit_buffer[15] ),
    .B(\soc/cpu/_02357_ ),
    .Y(\soc/cpu/_02361_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06746_  (.A1(\soc/cpu/_02360_ ),
    .A2(\soc/cpu/_02357_ ),
    .B1(\soc/cpu/_02361_ ),
    .Y(\soc/cpu/_00097_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_06747_  (.A_N(\soc/cpu/trap ),
    .B(_074_),
    .Y(\soc/cpu/_02362_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_06748_  (.A(\soc/cpu/mem_state[0] ),
    .B(\soc/cpu/mem_state[1] ),
    .Y(\soc/cpu/_02363_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06749_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_02362_ ),
    .C(\soc/cpu/_02363_ ),
    .Y(\soc/cpu/_02364_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_06750_  (.A(\soc/cpu/mem_state[0] ),
    .B(\soc/cpu/mem_state[1] ),
    .C(\soc/cpu/mem_do_wdata ),
    .D(\soc/cpu/_02362_ ),
    .X(\soc/cpu/_02365_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06751_  (.A(\soc/cpu/mem_do_rdata ),
    .B(\soc/cpu/_00711_ ),
    .C(\soc/cpu/_02365_ ),
    .Y(\soc/cpu/_02366_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06752_  (.A(\soc/cpu/mem_state[0] ),
    .B(\soc/cpu/mem_state[1] ),
    .Y(\soc/cpu/_02367_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06754_  (.A(_074_),
    .B(\soc/cpu/trap ),
    .Y(\soc/cpu/_02369_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06755_  (.A1(\soc/cpu/_02367_ ),
    .A2(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02369_ ),
    .B2(\soc/mem_ready ),
    .Y(\soc/cpu/_02370_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06756_  (.A(\soc/cpu/_02364_ ),
    .B(\soc/cpu/_02366_ ),
    .C(\soc/cpu/_02370_ ),
    .Y(\soc/cpu/_02371_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06757_  (.A_N(\soc/cpu/mem_do_wdata ),
    .B(\soc/cpu/_00715_ ),
    .Y(\soc/cpu/_02372_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06758_  (.A(\soc/cpu/_00745_ ),
    .B(\soc/cpu/_02350_ ),
    .Y(\soc/cpu/_02373_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06759_  (.A1(\soc/cpu/_02363_ ),
    .A2(\soc/cpu/_02372_ ),
    .B1(\soc/cpu/_02373_ ),
    .Y(\soc/cpu/_02374_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06760_  (.A1(\soc/cpu/_02362_ ),
    .A2(\soc/cpu/_02374_ ),
    .B1(\soc/cpu/_02371_ ),
    .Y(\soc/cpu/_02375_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_06761_  (.A1(\soc/mem_valid ),
    .A2(\soc/cpu/_02371_ ),
    .B1(\soc/cpu/_02375_ ),
    .X(\soc/cpu/_00098_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06762_  (.A(\soc/cpu/mem_la_read ),
    .B(\soc/cpu/_00857_ ),
    .Y(\soc/cpu/_02376_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06763_  (.A1(\soc/cpu/_00857_ ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_02376_ ),
    .B2(\iomem_wstrb[0] ),
    .X(\soc/cpu/_02377_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_06764_  (.A(\soc/cpu/_00743_ ),
    .B(\soc/cpu/_02352_ ),
    .X(\soc/cpu/_02378_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06765_  (.A1(\iomem_wstrb[0] ),
    .A2(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02377_ ),
    .B2(\soc/cpu/_02378_ ),
    .X(\soc/cpu/_00101_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06766_  (.A1(\soc/cpu/_00857_ ),
    .A2(\soc/cpu/mem_la_wstrb [1]),
    .B1(\soc/cpu/_02376_ ),
    .B2(\iomem_wstrb[1] ),
    .X(\soc/cpu/_02379_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06767_  (.A1(\iomem_wstrb[1] ),
    .A2(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02378_ ),
    .B2(\soc/cpu/_02379_ ),
    .X(\soc/cpu/_00102_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06768_  (.A1(\soc/cpu/_00857_ ),
    .A2(\soc/cpu/mem_la_wstrb [2]),
    .B1(\soc/cpu/_02376_ ),
    .B2(net404),
    .X(\soc/cpu/_02380_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06769_  (.A1(net404),
    .A2(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02378_ ),
    .B2(\soc/cpu/_02380_ ),
    .X(\soc/cpu/_00103_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06770_  (.A1(\soc/cpu/_00857_ ),
    .A2(\soc/cpu/mem_la_wstrb [3]),
    .B1(\soc/cpu/_02376_ ),
    .B2(\iomem_wstrb[3] ),
    .X(\soc/cpu/_02381_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06771_  (.A1(\iomem_wstrb[3] ),
    .A2(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02378_ ),
    .B2(\soc/cpu/_02381_ ),
    .X(\soc/cpu/_00104_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_06772_  (.A(\soc/cpu/mem_do_wdata ),
    .B(\soc/cpu/_00742_ ),
    .C(\soc/cpu/_02352_ ),
    .Y(\soc/cpu/_02382_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_06774_  (.A1(\soc/cpu/_00743_ ),
    .A2(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02382_ ),
    .C1(\soc/mem_instr ),
    .Y(\soc/cpu/_02384_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06775_  (.A1(\soc/cpu/_01159_ ),
    .A2(\soc/cpu/_02365_ ),
    .B1(\soc/cpu/_02384_ ),
    .Y(\soc/cpu/_00105_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_06777_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01110_ ),
    .C(\soc/cpu/_01116_ ),
    .Y(\soc/cpu/_02386_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_06778_  (.A(\soc/cpu/_01088_ ),
    .B(\soc/cpu/_01289_ ),
    .C(\soc/cpu/_01102_ ),
    .Y(\soc/cpu/_02387_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_06779_  (.A(\soc/cpu/_01363_ ),
    .B(\soc/cpu/_01124_ ),
    .C(\soc/cpu/_01233_ ),
    .D(\soc/cpu/_01272_ ),
    .Y(\soc/cpu/_02388_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06780_  (.A(\soc/cpu/_01189_ ),
    .B(\soc/cpu/_01363_ ),
    .C(\soc/cpu/_01117_ ),
    .Y(\soc/cpu/_02389_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_06781_  (.A1(\soc/cpu/_02386_ ),
    .A2(\soc/cpu/_02387_ ),
    .B1(\soc/cpu/_02388_ ),
    .C1(\soc/cpu/_02389_ ),
    .Y(\soc/cpu/_02390_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06783_  (.A(\soc/cpu/is_alu_reg_reg ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02392_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06784_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02390_ ),
    .B1(\soc/cpu/_02392_ ),
    .Y(\soc/cpu/_00106_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06785_  (.A(\soc/cpu/_01088_ ),
    .B(\soc/cpu/_01095_ ),
    .Y(\soc/cpu/_02393_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06786_  (.A(\soc/cpu/_02393_ ),
    .B(\soc/cpu/_01102_ ),
    .Y(\soc/cpu/_02394_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06787_  (.A(\soc/cpu/_02386_ ),
    .B(\soc/cpu/_02394_ ),
    .Y(\soc/cpu/_02395_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06788_  (.A(\soc/cpu/_01117_ ),
    .B(\soc/cpu/_01215_ ),
    .Y(\soc/cpu/_02396_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06789_  (.A(\soc/cpu/_01327_ ),
    .B(\soc/cpu/_02396_ ),
    .Y(\soc/cpu/_02397_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06790_  (.A(\soc/cpu/_01173_ ),
    .B(\soc/cpu/_02397_ ),
    .Y(\soc/cpu/_02398_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06791_  (.A(\soc/cpu/_01215_ ),
    .B(\soc/cpu/_01171_ ),
    .Y(\soc/cpu/_02399_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06792_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01164_ ),
    .Y(\soc/cpu/_02400_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06793_  (.A1(\soc/cpu/_01362_ ),
    .A2(\soc/cpu/_02399_ ),
    .B1(\soc/cpu/_02400_ ),
    .Y(\soc/cpu/_02401_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_06794_  (.A(\soc/cpu/_01183_ ),
    .B(\soc/cpu/_02398_ ),
    .C(\soc/cpu/_02401_ ),
    .X(\soc/cpu/_02402_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06795_  (.A(\soc/cpu/_02393_ ),
    .B(\soc/cpu/_01154_ ),
    .C(\soc/cpu/_02399_ ),
    .Y(\soc/cpu/_02403_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06796_  (.A(\soc/cpu/_01215_ ),
    .B(\soc/cpu/_01236_ ),
    .Y(\soc/cpu/_02404_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_06797_  (.A1(\soc/cpu/_01237_ ),
    .A2(\soc/cpu/_02403_ ),
    .B1(\soc/cpu/_02404_ ),
    .B2(\soc/cpu/_01189_ ),
    .Y(\soc/cpu/_02405_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06798_  (.A1(\soc/cpu/_01367_ ),
    .A2(\soc/cpu/_02402_ ),
    .B1(\soc/cpu/_02405_ ),
    .Y(\soc/cpu/_02406_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06799_  (.A(\soc/cpu/is_alu_reg_imm ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02407_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06800_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02395_ ),
    .A3(\soc/cpu/_02406_ ),
    .B1(\soc/cpu/_02407_ ),
    .Y(\soc/cpu/_00107_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_06801_  (.A_N(\soc/cpu/decoder_pseudo_trigger ),
    .B(\soc/cpu/decoder_trigger ),
    .Y(\soc/cpu/_02408_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_06804_  (.A(\soc/cpu/_00746_ ),
    .B(net784),
    .Y(\soc/cpu/_02411_ ));
 sky130_fd_sc_hd__and2_4 \soc/cpu/_06805_  (.A(net697),
    .B(\soc/cpu/_02411_ ),
    .X(\soc/cpu/_02412_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_06808_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .SLEEP(net951),
    .X(\soc/cpu/_02415_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06809_  (.A(\soc/cpu/mem_rdata_q[26] ),
    .B(\soc/cpu/mem_rdata_q[27] ),
    .Y(\soc/cpu/_02416_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06810_  (.A(\soc/cpu/mem_rdata_q[28] ),
    .B(\soc/cpu/mem_rdata_q[25] ),
    .Y(\soc/cpu/_02417_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06811_  (.A(\soc/cpu/mem_rdata_q[29] ),
    .B(\soc/cpu/mem_rdata_q[30] ),
    .C(\soc/cpu/mem_rdata_q[31] ),
    .Y(\soc/cpu/_02418_ ));
 sky130_fd_sc_hd__and3_4 \soc/cpu/_06812_  (.A(\soc/cpu/_02416_ ),
    .B(\soc/cpu/_02417_ ),
    .C(\soc/cpu/_02418_ ),
    .X(\soc/cpu/_02419_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06813_  (.A(\soc/cpu/_02415_ ),
    .B(\soc/cpu/_02419_ ),
    .Y(\soc/cpu/_02420_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06814_  (.A(\soc/cpu/_02416_ ),
    .B(\soc/cpu/_02417_ ),
    .Y(\soc/cpu/_02421_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06815_  (.A_N(\soc/cpu/mem_rdata_q[29] ),
    .B(\soc/cpu/mem_rdata_q[30] ),
    .Y(\soc/cpu/_02422_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_06816_  (.A(\soc/cpu/mem_rdata_q[31] ),
    .B(\soc/cpu/_02421_ ),
    .C(\soc/cpu/_02422_ ),
    .Y(\soc/cpu/_02423_ ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_06817_  (.A(net950),
    .B(\soc/cpu/_02415_ ),
    .X(\soc/cpu/_02424_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06818_  (.A(\soc/cpu/_02423_ ),
    .B(\soc/cpu/_02424_ ),
    .Y(\soc/cpu/_02425_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06819_  (.A(\soc/cpu/_02420_ ),
    .B(\soc/cpu/_02425_ ),
    .Y(\soc/cpu/_02426_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_06820_  (.A1(\soc/cpu/is_slli_srli_srai ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_02426_ ),
    .X(\soc/cpu/_00109_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_06821_  (.A(\soc/cpu/mem_rdata_q[27] ),
    .B(\soc/cpu/mem_rdata_q[29] ),
    .C(\soc/cpu/mem_rdata_q[30] ),
    .D(\soc/cpu/mem_rdata_q[31] ),
    .Y(\soc/cpu/_02427_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06822_  (.A(\soc/cpu/mem_rdata_q[25] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02428_ ));
 sky130_fd_sc_hd__nand3b_2 \soc/cpu/_06823_  (.A_N(\soc/cpu/mem_rdata_q[2] ),
    .B(\soc/cpu/mem_rdata_q[1] ),
    .C(\soc/cpu/mem_rdata_q[0] ),
    .Y(\soc/cpu/_02429_ ));
 sky130_fd_sc_hd__or4b_2 \soc/cpu/_06824_  (.A(\soc/cpu/mem_rdata_q[6] ),
    .B(\soc/cpu/mem_rdata_q[4] ),
    .C(\soc/cpu/mem_rdata_q[5] ),
    .D_N(\soc/cpu/mem_rdata_q[3] ),
    .X(\soc/cpu/_02430_ ));
 sky130_fd_sc_hd__nor4_4 \soc/cpu/_06825_  (.A(\soc/cpu/mem_rdata_q[28] ),
    .B(\soc/cpu/_02428_ ),
    .C(\soc/cpu/_02429_ ),
    .D(\soc/cpu/_02430_ ),
    .Y(\soc/cpu/_02431_ ));
 sky130_fd_sc_hd__a32o_1 \soc/cpu/_06829_  (.A1(\soc/cpu/mem_rdata_q[26] ),
    .A2(\soc/cpu/_02427_ ),
    .A3(\soc/cpu/_02431_ ),
    .B1(\soc/cpu/_02408_ ),
    .B2(\soc/cpu/instr_maskirq ),
    .X(\soc/cpu/_00110_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06830_  (.A(\soc/cpu/_01088_ ),
    .B(\soc/cpu/_01095_ ),
    .C(\soc/cpu/_01102_ ),
    .X(\soc/cpu/_02435_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06831_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01110_ ),
    .C(\soc/cpu/_01241_ ),
    .Y(\soc/cpu/_02436_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06832_  (.A(\soc/cpu/_02435_ ),
    .B(\soc/cpu/_02436_ ),
    .Y(\soc/cpu/_02437_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06833_  (.A(\soc/cpu/_01258_ ),
    .B(\soc/cpu/_01270_ ),
    .C(\soc/cpu/_01590_ ),
    .Y(\soc/cpu/_02438_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06834_  (.A(\soc/cpu/_01053_ ),
    .B(\soc/cpu/_01246_ ),
    .Y(\soc/cpu/_02439_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06835_  (.A(\soc/cpu/_02438_ ),
    .B(\soc/cpu/_02439_ ),
    .Y(\soc/cpu/_02440_ ));
 sky130_fd_sc_hd__or4_4 \soc/cpu/_06836_  (.A(\soc/cpu/_01205_ ),
    .B(\soc/cpu/_01224_ ),
    .C(\soc/cpu/_02437_ ),
    .D(\soc/cpu/_02440_ ),
    .X(\soc/cpu/_02441_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06838_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02443_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06839_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02441_ ),
    .B1(\soc/cpu/_02443_ ),
    .Y(\soc/cpu/_00111_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06840_  (.A(\soc/cpu/decoded_imm_j[1] ),
    .Y(\soc/cpu/_02444_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_06841_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02445_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_06842_  (.A(\soc/cpu/mem_do_rinst ),
    .B(\soc/cpu/_00963_ ),
    .Y(\soc/cpu/_02446_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_06844_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02448_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06845_  (.A(\soc/cpu/_01369_ ),
    .B(\soc/cpu/_02448_ ),
    .Y(\soc/cpu/_02449_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/_06846_  (.A1(\soc/cpu/_02444_ ),
    .A2(\soc/cpu/_01588_ ),
    .B1(\soc/cpu/_02445_ ),
    .B2(\soc/cpu/_01241_ ),
    .C1(\soc/cpu/_02449_ ),
    .Y(\soc/cpu/_00112_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06847_  (.A(\soc/cpu/_01376_ ),
    .B(\soc/cpu/_02448_ ),
    .Y(\soc/cpu/_02450_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06849_  (.A(\soc/cpu/_01102_ ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02452_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06850_  (.A1(\soc/cpu/decoded_imm_j[2] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02452_ ),
    .B2(\soc/cpu/_00738_ ),
    .Y(\soc/cpu/_02453_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06851_  (.A(\soc/cpu/_02450_ ),
    .B(\soc/cpu/_02453_ ),
    .Y(\soc/cpu/_00113_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06852_  (.A(\soc/cpu/decoded_imm_j[3] ),
    .Y(\soc/cpu/_02454_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06854_  (.A(\soc/cpu/_00730_ ),
    .B(\soc/cpu/_00737_ ),
    .C(\soc/cpu/_01386_ ),
    .X(\soc/cpu/_02456_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_06855_  (.A1(\soc/cpu/_00738_ ),
    .A2(\soc/cpu/_01210_ ),
    .B1(\soc/cpu/_02446_ ),
    .C1(\soc/cpu/_02456_ ),
    .Y(\soc/cpu/_02457_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06856_  (.A1(\soc/cpu/_02454_ ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02457_ ),
    .Y(\soc/cpu/_00114_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06857_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01396_ ),
    .Y(\soc/cpu/_02458_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06858_  (.A(\soc/cpu/decoded_imm_j[4] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02459_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06859_  (.A1(\soc/cpu/_01300_ ),
    .A2(\soc/cpu/_01588_ ),
    .A3(\soc/cpu/_02458_ ),
    .B1(\soc/cpu/_02459_ ),
    .Y(\soc/cpu/_00115_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06861_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02461_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_06862_  (.A1(\soc/cpu/decoded_imm_j[5] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02461_ ),
    .B2(\soc/cpu/_01110_ ),
    .C1(\soc/cpu/_02448_ ),
    .C2(\soc/cpu/_01053_ ),
    .Y(\soc/cpu/_02462_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06863_  (.A(\soc/cpu/_02462_ ),
    .Y(\soc/cpu/_00116_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_06864_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02463_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06865_  (.A(\soc/cpu/decoded_imm_j[6] ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02464_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/_06866_  (.A1(\soc/cpu/_01146_ ),
    .A2(\soc/cpu/_02445_ ),
    .B1(\soc/cpu/_02463_ ),
    .B2(\soc/cpu/_01205_ ),
    .C1(\soc/cpu/_02464_ ),
    .Y(\soc/cpu/_00117_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06867_  (.A1(\soc/cpu/decoded_imm_j[7] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02448_ ),
    .B2(\soc/cpu/_01224_ ),
    .Y(\soc/cpu/_02465_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06868_  (.A1(\soc/cpu/_01095_ ),
    .A2(\soc/cpu/_02445_ ),
    .B1(\soc/cpu/_02465_ ),
    .Y(\soc/cpu/_00118_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06869_  (.A1(\soc/cpu/decoded_imm_j[8] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02448_ ),
    .B2(\soc/cpu/_01246_ ),
    .Y(\soc/cpu/_02466_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06870_  (.A1(\soc/cpu/_01140_ ),
    .A2(\soc/cpu/_02445_ ),
    .B1(\soc/cpu/_02466_ ),
    .Y(\soc/cpu/_00119_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06871_  (.A1(\soc/cpu/decoded_imm_j[9] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02448_ ),
    .B2(\soc/cpu/_01258_ ),
    .Y(\soc/cpu/_02467_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06872_  (.A1(\soc/cpu/_01152_ ),
    .A2(\soc/cpu/_02445_ ),
    .B1(\soc/cpu/_02467_ ),
    .Y(\soc/cpu/_00120_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_06873_  (.A1(\soc/cpu/decoded_imm_j[10] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02461_ ),
    .B2(\soc/cpu/_01137_ ),
    .C1(\soc/cpu/_02448_ ),
    .C2(\soc/cpu/_01270_ ),
    .Y(\soc/cpu/_02468_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06874_  (.A(\soc/cpu/_02468_ ),
    .Y(\soc/cpu/_00121_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06875_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01124_ ),
    .Y(\soc/cpu/_02469_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06876_  (.A1(\soc/cpu/_00827_ ),
    .A2(\soc/cpu/_01356_ ),
    .B1(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02470_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06877_  (.A(\soc/cpu/decoded_imm_j[11] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02471_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06878_  (.A1(\soc/cpu/_02469_ ),
    .A2(\soc/cpu/_02470_ ),
    .B1(\soc/cpu/_02471_ ),
    .Y(\soc/cpu/_00122_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06880_  (.A(\soc/cpu/decoded_imm_j[12] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02473_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06881_  (.A1(\soc/cpu/_01215_ ),
    .A2(\soc/cpu/_01588_ ),
    .B1(\soc/cpu/_02473_ ),
    .Y(\soc/cpu/_00123_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_06882_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01215_ ),
    .C(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02474_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06883_  (.A1(\soc/cpu/decoded_imm_j[13] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02474_ ),
    .Y(\soc/cpu/_02475_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06884_  (.A1(\soc/cpu/_01072_ ),
    .A2(\soc/cpu/_02463_ ),
    .B1(\soc/cpu/_02475_ ),
    .Y(\soc/cpu/_00124_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06885_  (.A1(\soc/cpu/decoded_imm_j[14] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02474_ ),
    .Y(\soc/cpu/_02476_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06886_  (.A1(\soc/cpu/_01164_ ),
    .A2(\soc/cpu/_02463_ ),
    .B1(\soc/cpu/_02476_ ),
    .Y(\soc/cpu/_00125_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06887_  (.A1(\soc/cpu/decoded_imm_j[15] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02474_ ),
    .Y(\soc/cpu/_02477_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06888_  (.A1(\soc/cpu/_01169_ ),
    .A2(\soc/cpu/_02463_ ),
    .B1(\soc/cpu/_02477_ ),
    .Y(\soc/cpu/_00126_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06889_  (.A1(\soc/cpu/decoded_imm_j[16] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02474_ ),
    .Y(\soc/cpu/_02478_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06890_  (.A1(\soc/cpu/_01342_ ),
    .A2(\soc/cpu/_02463_ ),
    .B1(\soc/cpu/_02478_ ),
    .Y(\soc/cpu/_00127_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06891_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01124_ ),
    .C(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02479_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06892_  (.A(\soc/cpu/_01345_ ),
    .B(\soc/cpu/_02463_ ),
    .Y(\soc/cpu/_02480_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06893_  (.A1(\soc/cpu/decoded_imm_j[17] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02480_ ),
    .Y(\soc/cpu/_02481_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06894_  (.A(\soc/cpu/_02479_ ),
    .B(\soc/cpu/_02481_ ),
    .Y(\soc/cpu/_00128_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06895_  (.A1(\soc/cpu/decoded_imm_j[18] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02474_ ),
    .Y(\soc/cpu/_02482_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06896_  (.A1(\soc/cpu/_01351_ ),
    .A2(\soc/cpu/_02463_ ),
    .B1(\soc/cpu/_02482_ ),
    .Y(\soc/cpu/_00129_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06897_  (.A1(\soc/cpu/decoded_imm_j[19] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02448_ ),
    .B2(\soc/cpu/_01354_ ),
    .Y(\soc/cpu/_02483_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06898_  (.A(\soc/cpu/_02479_ ),
    .B(\soc/cpu/_02483_ ),
    .Y(\soc/cpu/_00130_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_06899_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .Y(\soc/cpu/_02484_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06900_  (.A1(\soc/cpu/_01590_ ),
    .A2(\soc/cpu/_02448_ ),
    .B1(\soc/cpu/_02474_ ),
    .Y(\soc/cpu/_02485_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06901_  (.A1(\soc/cpu/_02484_ ),
    .A2(\soc/cpu/_01588_ ),
    .B1(\soc/cpu/_02485_ ),
    .Y(\soc/cpu/_00131_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_06902_  (.A(\soc/cpu/mem_rdata_q[27] ),
    .SLEEP(\soc/cpu/mem_rdata_q[26] ),
    .X(\soc/cpu/_02486_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06903_  (.A(\soc/cpu/mem_rdata_q[25] ),
    .B(\soc/cpu/mem_rdata_q[24] ),
    .Y(\soc/cpu/_02487_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06904_  (.A(\soc/cpu/_02486_ ),
    .B(\soc/cpu/_02487_ ),
    .Y(\soc/cpu/_02488_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06905_  (.A(\soc/cpu/mem_rdata_q[22] ),
    .B(\soc/cpu/mem_rdata_q[20] ),
    .C(\soc/cpu/mem_rdata_q[23] ),
    .Y(\soc/cpu/_02489_ ));
 sky130_fd_sc_hd__nor4b_1 \soc/cpu/_06906_  (.A(\soc/cpu/mem_rdata_q[3] ),
    .B(\soc/cpu/_02422_ ),
    .C(\soc/cpu/mem_rdata_q[28] ),
    .D_N(\soc/cpu/mem_rdata_q[31] ),
    .Y(\soc/cpu/_02490_ ));
 sky130_fd_sc_hd__or3b_4 \soc/cpu/_06907_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(net950),
    .C_N(net951),
    .X(\soc/cpu/_02491_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06908_  (.A(\soc/cpu/mem_rdata_q[19] ),
    .B(\soc/cpu/_02491_ ),
    .Y(\soc/cpu/_02492_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06909_  (.A(\soc/cpu/mem_rdata_q[6] ),
    .B(\soc/cpu/mem_rdata_q[4] ),
    .C(\soc/cpu/mem_rdata_q[5] ),
    .Y(\soc/cpu/_02493_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_06910_  (.A(\soc/cpu/mem_rdata_q[16] ),
    .B(\soc/cpu/mem_rdata_q[17] ),
    .C(\soc/cpu/mem_rdata_q[18] ),
    .D(\soc/cpu/mem_rdata_q[15] ),
    .X(\soc/cpu/_02494_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_06911_  (.A(\soc/cpu/_02408_ ),
    .B(\soc/cpu/_02429_ ),
    .C(\soc/cpu/_02493_ ),
    .D(\soc/cpu/_02494_ ),
    .Y(\soc/cpu/_02495_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/_06912_  (.A(\soc/cpu/_02490_ ),
    .B(\soc/cpu/_02492_ ),
    .C(\soc/cpu/_02495_ ),
    .Y(\soc/cpu/_02496_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_06913_  (.A(\soc/cpu/_02496_ ),
    .Y(\soc/cpu/_02497_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06914_  (.A(\soc/cpu/mem_rdata_q[21] ),
    .B(\soc/cpu/_02489_ ),
    .C(\soc/cpu/_02497_ ),
    .Y(\soc/cpu/_02498_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06916_  (.A(\soc/cpu/instr_rdinstrh ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02500_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06917_  (.A1(\soc/cpu/_02488_ ),
    .A2(\soc/cpu/_02498_ ),
    .B1(\soc/cpu/_02500_ ),
    .Y(\soc/cpu/_00132_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_06918_  (.A(\soc/cpu/mem_rdata_q[22] ),
    .B(\soc/cpu/mem_rdata_q[21] ),
    .C(\soc/cpu/mem_rdata_q[23] ),
    .X(\soc/cpu/_02501_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06920_  (.A(\soc/cpu/instr_rdcycleh ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02503_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06921_  (.A1(\soc/cpu/_02488_ ),
    .A2(\soc/cpu/_02496_ ),
    .A3(\soc/cpu/_02501_ ),
    .B1(\soc/cpu/_02503_ ),
    .Y(\soc/cpu/_00134_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06922_  (.A(\soc/cpu/_02416_ ),
    .B(\soc/cpu/_02487_ ),
    .Y(\soc/cpu/_02504_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06923_  (.A(\soc/cpu/instr_rdcycle ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02505_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_06924_  (.A1(\soc/cpu/_02496_ ),
    .A2(\soc/cpu/_02501_ ),
    .A3(\soc/cpu/_02504_ ),
    .B1(\soc/cpu/_02505_ ),
    .Y(\soc/cpu/_00135_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06925_  (.A(\soc/cpu/instr_srli ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02506_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06926_  (.A(\soc/cpu/_02412_ ),
    .B(\soc/cpu/_02419_ ),
    .C(\soc/cpu/_02424_ ),
    .Y(\soc/cpu/_02507_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06927_  (.A(\soc/cpu/_02506_ ),
    .B(\soc/cpu/_02507_ ),
    .Y(\soc/cpu/_00144_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_06928_  (.A_N(\soc/cpu/mem_rdata_q[13] ),
    .B(\soc/cpu/mem_rdata_q[12] ),
    .Y(\soc/cpu/_02508_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06929_  (.A(net950),
    .B(\soc/cpu/_02508_ ),
    .Y(\soc/cpu/_02509_ ));
 sky130_fd_sc_hd__a32o_1 \soc/cpu/_06930_  (.A1(\soc/cpu/_02412_ ),
    .A2(\soc/cpu/_02419_ ),
    .A3(\soc/cpu/_02509_ ),
    .B1(\soc/cpu/_02408_ ),
    .B2(\soc/cpu/instr_slli ),
    .X(\soc/cpu/_00145_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06932_  (.A(net952),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02511_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06934_  (.A(\soc/cpu/instr_sw ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02513_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06935_  (.A1(\soc/cpu/_02491_ ),
    .A2(\soc/cpu/_02511_ ),
    .B1(\soc/cpu/_02513_ ),
    .Y(\soc/cpu/_00146_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_06936_  (.A(net950),
    .B(\soc/cpu/_02508_ ),
    .X(\soc/cpu/_02514_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06937_  (.A(\soc/cpu/instr_sh ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02515_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06938_  (.A1(\soc/cpu/_02514_ ),
    .A2(\soc/cpu/_02511_ ),
    .B1(\soc/cpu/_02515_ ),
    .Y(\soc/cpu/_00153_ ));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_06939_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(net951),
    .C(net950),
    .X(\soc/cpu/_02516_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06940_  (.A(\soc/cpu/instr_sb ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02517_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06941_  (.A1(\soc/cpu/_02511_ ),
    .A2(\soc/cpu/_02516_ ),
    .B1(\soc/cpu/_02517_ ),
    .Y(\soc/cpu/_00154_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06942_  (.A(net852),
    .B(\soc/cpu/_02415_ ),
    .Y(\soc/cpu/_02518_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06943_  (.A(net953),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02519_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06944_  (.A(\soc/cpu/instr_lhu ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02520_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06945_  (.A1(\soc/cpu/_02518_ ),
    .A2(\soc/cpu/_02519_ ),
    .B1(\soc/cpu/_02520_ ),
    .Y(\soc/cpu/_00155_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06946_  (.A(\soc/cpu/instr_lbu ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02521_ ));
 sky130_fd_sc_hd__nor3b_2 \soc/cpu/_06948_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(net951),
    .C_N(net950),
    .Y(\soc/cpu/_02523_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06949_  (.A(net953),
    .B(\soc/cpu/_02411_ ),
    .C(\soc/cpu/_02523_ ),
    .Y(\soc/cpu/_02524_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06950_  (.A(\soc/cpu/_02521_ ),
    .B(\soc/cpu/_02524_ ),
    .Y(\soc/cpu/_00156_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06951_  (.A(\soc/cpu/instr_lh ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02525_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06952_  (.A1(\soc/cpu/_02514_ ),
    .A2(\soc/cpu/_02519_ ),
    .B1(\soc/cpu/_02525_ ),
    .Y(\soc/cpu/_00157_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06953_  (.A(\soc/cpu/_02400_ ),
    .B(\soc/cpu/_01124_ ),
    .Y(\soc/cpu/_02526_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06954_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01110_ ),
    .C(\soc/cpu/_01241_ ),
    .X(\soc/cpu/_02527_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_06955_  (.A(\soc/cpu/_01210_ ),
    .B(\soc/cpu/_01289_ ),
    .C(\soc/cpu/_01102_ ),
    .X(\soc/cpu/_02528_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_06956_  (.A(\soc/cpu/_01189_ ),
    .B(\soc/cpu/_01118_ ),
    .C(\soc/cpu/_01155_ ),
    .Y(\soc/cpu/_02529_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06957_  (.A1(\soc/cpu/_02526_ ),
    .A2(\soc/cpu/_02527_ ),
    .A3(\soc/cpu/_02528_ ),
    .B1(\soc/cpu/_02529_ ),
    .Y(\soc/cpu/_02530_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06958_  (.A(\soc/cpu/instr_jalr ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02531_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06959_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02530_ ),
    .B1(\soc/cpu/_02531_ ),
    .Y(\soc/cpu/_00158_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_06960_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01110_ ),
    .C(\soc/cpu/_01116_ ),
    .D(\soc/cpu/_02528_ ),
    .Y(\soc/cpu/_02532_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06963_  (.A(\soc/cpu/instr_jal ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02535_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_06964_  (.A1(\soc/cpu/_01248_ ),
    .A2(\soc/cpu/_01588_ ),
    .A3(\soc/cpu/_02532_ ),
    .B1(\soc/cpu/_02535_ ),
    .Y(\soc/cpu/_00163_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_06965_  (.A(\soc/cpu/_02394_ ),
    .B(\soc/cpu/_02527_ ),
    .Y(\soc/cpu/_02536_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06966_  (.A(\soc/cpu/instr_auipc ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02537_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06967_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02536_ ),
    .B1(\soc/cpu/_02537_ ),
    .Y(\soc/cpu/_00164_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_06968_  (.A0(\soc/cpu/latched_compr ),
    .A1(\soc/cpu/compressed_instr ),
    .S(\soc/cpu/_00796_ ),
    .X(\soc/cpu/_00166_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06969_  (.A(\soc/cpu/cpuregs_rdata2[0] ),
    .B(\soc/cpu/_00957_ ),
    .C(\soc/cpu/_01414_ ),
    .Y(\soc/cpu/_02538_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06971_  (.A1(\soc/cpu/decoded_imm[0] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02540_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06973_  (.A(\soc/cpu/mem_la_wdata [0]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02542_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06974_  (.A1(\soc/cpu/_02538_ ),
    .A2(\soc/cpu/_02540_ ),
    .B1(\soc/cpu/_02542_ ),
    .Y(\soc/cpu/_00247_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06976_  (.A(\soc/cpu/cpuregs_rdata2[1] ),
    .B(\soc/cpu/_00957_ ),
    .C(\soc/cpu/_01414_ ),
    .Y(\soc/cpu/_02544_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06978_  (.A1(\soc/cpu/decoded_imm[1] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02546_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06979_  (.A1(\soc/cpu/_01521_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02544_ ),
    .B2(\soc/cpu/_02546_ ),
    .Y(\soc/cpu/_00248_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06980_  (.A(\soc/cpu/cpuregs_rdata2[2] ),
    .B(\soc/cpu/_00957_ ),
    .C(\soc/cpu/_01414_ ),
    .Y(\soc/cpu/_02547_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06981_  (.A1(\soc/cpu/decoded_imm[2] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02548_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06982_  (.A1(\soc/cpu/_01520_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02547_ ),
    .B2(\soc/cpu/_02548_ ),
    .Y(\soc/cpu/_00249_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_06983_  (.A(\soc/cpu/cpuregs_rdata2[3] ),
    .B(\soc/cpu/_00957_ ),
    .C(\soc/cpu/_01414_ ),
    .Y(\soc/cpu/_02549_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06984_  (.A1(net857),
    .A2(\soc/cpu/_00966_ ),
    .B1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02550_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_06985_  (.A1(\soc/cpu/_01519_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02549_ ),
    .B2(\soc/cpu/_02550_ ),
    .Y(\soc/cpu/_00250_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_06987_  (.A1(\soc/cpu/_00966_ ),
    .A2(\soc/cpu/_01426_ ),
    .B1(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02552_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06988_  (.A1(\soc/cpu/decoded_imm[4] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(\soc/cpu/_02552_ ),
    .Y(\soc/cpu/_02553_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06989_  (.A1(\soc/cpu/_01518_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02553_ ),
    .Y(\soc/cpu/_00251_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_06990_  (.A1(\soc/cpu/_01412_ ),
    .A2(\soc/cpu/_01413_ ),
    .B1(\soc/cpu/_00966_ ),
    .Y(\soc/cpu/_02554_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_06993_  (.A1(\soc/cpu/decoded_imm[5] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[5] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02557_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_06994_  (.A1(\soc/cpu/_01517_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02557_ ),
    .Y(\soc/cpu/_00252_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06995_  (.A(\soc/cpu/mem_la_wdata [6]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02558_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_06997_  (.A1(\soc/cpu/decoded_imm[6] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[6] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02560_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_06998_  (.A(\soc/cpu/_02558_ ),
    .B(\soc/cpu/_02560_ ),
    .Y(\soc/cpu/_00253_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_06999_  (.A1(\soc/cpu/decoded_imm[7] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[7] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02561_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07000_  (.A1(\soc/cpu/_01516_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02561_ ),
    .Y(\soc/cpu/_00254_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07001_  (.A(\soc/cpu/pcpi_rs2 [8]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02562_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07002_  (.A1(\soc/cpu/decoded_imm[8] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[8] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02563_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07003_  (.A(\soc/cpu/_02562_ ),
    .B(\soc/cpu/_02563_ ),
    .Y(\soc/cpu/_00255_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07004_  (.A1(\soc/cpu/decoded_imm[9] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[9] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02564_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07005_  (.A1(\soc/cpu/_01538_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02564_ ),
    .Y(\soc/cpu/_00256_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07006_  (.A1(net872),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[10] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02565_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07007_  (.A1(\soc/cpu/_01869_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02565_ ),
    .Y(\soc/cpu/_00257_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07008_  (.A1(\soc/cpu/decoded_imm[11] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[11] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02566_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07009_  (.A1(\soc/cpu/_01537_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02566_ ),
    .Y(\soc/cpu/_00258_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07011_  (.A1(net879),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[12] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02568_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07012_  (.A1(\soc/cpu/_01534_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02568_ ),
    .Y(\soc/cpu/_00259_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07013_  (.A1(\soc/cpu/decoded_imm[13] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[13] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02569_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07014_  (.A1(\soc/cpu/_01533_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02569_ ),
    .Y(\soc/cpu/_00260_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07015_  (.A(\soc/cpu/pcpi_rs2 [14]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02570_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07016_  (.A1(\soc/cpu/decoded_imm[14] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[14] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02571_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07017_  (.A(\soc/cpu/_02570_ ),
    .B(\soc/cpu/_02571_ ),
    .Y(\soc/cpu/_00261_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07018_  (.A1(\soc/cpu/decoded_imm[15] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[15] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02572_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07019_  (.A1(\soc/cpu/_01530_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02572_ ),
    .Y(\soc/cpu/_00262_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07020_  (.A(\soc/cpu/pcpi_rs2 [16]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02573_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07021_  (.A1(\soc/cpu/decoded_imm[16] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[16] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02574_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07022_  (.A(\soc/cpu/_02573_ ),
    .B(\soc/cpu/_02574_ ),
    .Y(\soc/cpu/_00263_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07023_  (.A(\soc/cpu/pcpi_rs2 [17]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02575_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07024_  (.A1(\soc/cpu/decoded_imm[17] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net144),
    .B2(\soc/cpu/cpuregs_rdata2[17] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02576_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07025_  (.A(\soc/cpu/_02575_ ),
    .B(\soc/cpu/_02576_ ),
    .Y(\soc/cpu/_00264_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07026_  (.A(\soc/cpu/pcpi_rs2 [18]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02577_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07027_  (.A1(\soc/cpu/decoded_imm[18] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(\soc/cpu/_02554_ ),
    .B2(\soc/cpu/cpuregs_rdata2[18] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02578_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07028_  (.A(\soc/cpu/_02577_ ),
    .B(\soc/cpu/_02578_ ),
    .Y(\soc/cpu/_00265_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07029_  (.A1(net890),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[19] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02579_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07030_  (.A1(\soc/cpu/_01554_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02579_ ),
    .Y(\soc/cpu/_00266_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07031_  (.A(\soc/cpu/pcpi_rs2 [20]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02580_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07032_  (.A1(net889),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[20] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02581_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07033_  (.A(\soc/cpu/_02580_ ),
    .B(\soc/cpu/_02581_ ),
    .Y(\soc/cpu/_00267_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07034_  (.A1(\soc/cpu/decoded_imm[21] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[21] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02582_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07035_  (.A1(\soc/cpu/_01551_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02582_ ),
    .Y(\soc/cpu/_00268_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07036_  (.A(\soc/cpu/pcpi_rs2 [22]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02583_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07037_  (.A1(\soc/cpu/decoded_imm[22] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[22] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02584_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07038_  (.A(\soc/cpu/_02583_ ),
    .B(\soc/cpu/_02584_ ),
    .Y(\soc/cpu/_00269_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07039_  (.A(\soc/cpu/pcpi_rs2 [23]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02585_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07040_  (.A1(\soc/cpu/decoded_imm[23] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[23] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02586_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07041_  (.A(\soc/cpu/_02585_ ),
    .B(\soc/cpu/_02586_ ),
    .Y(\soc/cpu/_00270_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07042_  (.A(\soc/cpu/pcpi_rs2 [24]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02587_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07043_  (.A1(\soc/cpu/decoded_imm[24] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[24] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02588_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07044_  (.A(\soc/cpu/_02587_ ),
    .B(\soc/cpu/_02588_ ),
    .Y(\soc/cpu/_00271_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07045_  (.A1(\soc/cpu/decoded_imm[25] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[25] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02589_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07046_  (.A1(\soc/cpu/_02037_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02589_ ),
    .Y(\soc/cpu/_00272_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07047_  (.A1(\soc/cpu/decoded_imm[26] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[26] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02590_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07048_  (.A1(\soc/cpu/_02053_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02590_ ),
    .Y(\soc/cpu/_00273_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07049_  (.A1(\soc/cpu/decoded_imm[27] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[27] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02591_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07050_  (.A1(\soc/cpu/_01569_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02591_ ),
    .Y(\soc/cpu/_00274_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07051_  (.A1(net854),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[28] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02592_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07052_  (.A1(\soc/cpu/_01568_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02592_ ),
    .Y(\soc/cpu/_00275_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07053_  (.A1(net853),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[29] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02593_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07054_  (.A1(\soc/cpu/_01567_ ),
    .A2(\soc/cpu/_00894_ ),
    .B1(\soc/cpu/_02593_ ),
    .Y(\soc/cpu/_00276_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07055_  (.A(\soc/cpu/pcpi_rs2 [30]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02594_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07056_  (.A1(\soc/cpu/decoded_imm[30] ),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[30] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02595_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07057_  (.A(\soc/cpu/_02594_ ),
    .B(\soc/cpu/_02595_ ),
    .Y(\soc/cpu/_00277_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07058_  (.A(\soc/cpu/pcpi_rs2 [31]),
    .B(\soc/cpu/_00906_ ),
    .Y(\soc/cpu/_02596_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07059_  (.A1(net878),
    .A2(\soc/cpu/_00966_ ),
    .B1(net143),
    .B2(\soc/cpu/cpuregs_rdata2[31] ),
    .C1(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_02597_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07060_  (.A(\soc/cpu/_02596_ ),
    .B(\soc/cpu/_02597_ ),
    .Y(\soc/cpu/_00278_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07061_  (.A(\soc/cpu/mem_do_wdata ),
    .B(\soc/cpu/cpu_state[5] ),
    .Y(\soc/cpu/_02598_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07062_  (.A1(\soc/cpu/_00842_ ),
    .A2(\soc/cpu/_02598_ ),
    .B1(\soc/cpu/_00838_ ),
    .Y(\soc/cpu/_02599_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07063_  (.A1(\soc/cpu/reg_sh[1] ),
    .A2(\soc/cpu/_00976_ ),
    .B1(\soc/cpu/cpu_state[4] ),
    .Y(\soc/cpu/_02600_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_07064_  (.A(\soc/cpu/instr_sra ),
    .B(\soc/cpu/instr_srai ),
    .Y(\soc/cpu/_02601_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07065_  (.A(\soc/cpu/instr_srl ),
    .B(\soc/cpu/instr_srli ),
    .Y(\soc/cpu/_02602_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_07066_  (.A(\soc/cpu/_02601_ ),
    .B(\soc/cpu/_02602_ ),
    .Y(\soc/cpu/_02603_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_07067_  (.A(\soc/cpu/instr_sll ),
    .B(\soc/cpu/instr_slli ),
    .C(\soc/cpu/_02600_ ),
    .D(\soc/cpu/_02603_ ),
    .X(\soc/cpu/_02604_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_07068_  (.A(_074_),
    .B(\soc/cpu/_00938_ ),
    .C(\soc/cpu/_00990_ ),
    .D(\soc/cpu/_02604_ ),
    .Y(\soc/cpu/_02605_ ));
 sky130_fd_sc_hd__a311oi_1 \soc/cpu/_07069_  (.A1(\soc/cpu/mem_do_rdata ),
    .A2(\soc/cpu/cpu_state[6] ),
    .A3(\soc/cpu/_00842_ ),
    .B1(\soc/cpu/_02599_ ),
    .C1(\soc/cpu/_02605_ ),
    .Y(\soc/cpu/_02606_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07071_  (.A1(\soc/cpu/instr_sra ),
    .A2(\soc/cpu/instr_srai ),
    .B1(\soc/cpu/_00979_ ),
    .Y(\soc/cpu/_02608_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07072_  (.A1(net47),
    .A2(\soc/cpu/_02608_ ),
    .B1(\soc/cpu/pcpi_rs1 [31]),
    .Y(\soc/cpu/_02609_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07073_  (.A(\soc/cpu/decoded_imm[30] ),
    .B(\soc/cpu/pcpi_rs1 [30]),
    .Y(\soc/cpu/_02610_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07074_  (.A(\soc/cpu/decoded_imm[29] ),
    .B(\soc/cpu/pcpi_rs1 [29]),
    .X(\soc/cpu/_02611_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07075_  (.A(\soc/cpu/decoded_imm[27] ),
    .B(\soc/cpu/pcpi_rs1 [27]),
    .Y(\soc/cpu/_02612_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07076_  (.A(\soc/cpu/decoded_imm[25] ),
    .B(\soc/cpu/pcpi_rs1 [25]),
    .Y(\soc/cpu/_02613_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07077_  (.A(\soc/cpu/decoded_imm[23] ),
    .B(\soc/cpu/pcpi_rs1 [23]),
    .Y(\soc/cpu/_02614_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_07078_  (.A(\soc/cpu/decoded_imm[22] ),
    .B(\soc/cpu/pcpi_rs1 [22]),
    .X(\soc/cpu/_02615_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07079_  (.A(\soc/cpu/decoded_imm[19] ),
    .B(\soc/cpu/pcpi_rs1 [19]),
    .Y(\soc/cpu/_02616_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07080_  (.A(\soc/cpu/decoded_imm[18] ),
    .B(\soc/cpu/pcpi_rs1 [18]),
    .X(\soc/cpu/_02617_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07081_  (.A(\soc/cpu/decoded_imm[18] ),
    .B(\soc/cpu/pcpi_rs1 [18]),
    .Y(\soc/cpu/_02618_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07082_  (.A(\soc/cpu/_02617_ ),
    .B(\soc/cpu/_02618_ ),
    .Y(\soc/cpu/_02619_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_07083_  (.A(\soc/cpu/decoded_imm[17] ),
    .B(\soc/cpu/pcpi_rs1 [17]),
    .X(\soc/cpu/_02620_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_07084_  (.A(\soc/cpu/decoded_imm[16] ),
    .B(\soc/cpu/pcpi_rs1 [16]),
    .Y(\soc/cpu/_02621_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07085_  (.A(\soc/cpu/decoded_imm[15] ),
    .B(\soc/cpu/pcpi_rs1 [15]),
    .Y(\soc/cpu/_02622_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_07086_  (.A(\soc/cpu/decoded_imm[14] ),
    .B(\soc/cpu/pcpi_rs1 [14]),
    .X(\soc/cpu/_02623_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07087_  (.A(\soc/cpu/decoded_imm[14] ),
    .B(\soc/cpu/pcpi_rs1 [14]),
    .Y(\soc/cpu/_02624_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07088_  (.A(\soc/cpu/_02623_ ),
    .B(\soc/cpu/_02624_ ),
    .Y(\soc/cpu/_02625_ ));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_07089_  (.A(\soc/cpu/decoded_imm[13] ),
    .B(\soc/cpu/pcpi_rs1 [13]),
    .X(\soc/cpu/_02626_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_07090_  (.A(\soc/cpu/decoded_imm[12] ),
    .B(\soc/cpu/pcpi_rs1 [12]),
    .Y(\soc/cpu/_02627_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07091_  (.A(\soc/cpu/decoded_imm[11] ),
    .B(\soc/cpu/pcpi_rs1 [11]),
    .Y(\soc/cpu/_02628_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_07092_  (.A(\soc/cpu/decoded_imm[10] ),
    .B(\soc/cpu/pcpi_rs1 [10]),
    .X(\soc/cpu/_02629_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07093_  (.A(\soc/cpu/decoded_imm[10] ),
    .B(\soc/cpu/pcpi_rs1 [10]),
    .Y(\soc/cpu/_02630_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07094_  (.A(\soc/cpu/_02629_ ),
    .B(\soc/cpu/_02630_ ),
    .Y(\soc/cpu/_02631_ ));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_07095_  (.A(\soc/cpu/decoded_imm[9] ),
    .B(\soc/cpu/pcpi_rs1 [9]),
    .X(\soc/cpu/_02632_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_07096_  (.A(\soc/cpu/decoded_imm[8] ),
    .B(\soc/cpu/pcpi_rs1 [8]),
    .Y(\soc/cpu/_02633_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07097_  (.A(\soc/cpu/decoded_imm[7] ),
    .B(\soc/cpu/pcpi_rs1 [7]),
    .Y(\soc/cpu/_02634_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07098_  (.A(\soc/cpu/decoded_imm[6] ),
    .B(\soc/cpu/pcpi_rs1 [6]),
    .Y(\soc/cpu/_02635_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07099_  (.A(\soc/cpu/decoded_imm[5] ),
    .B(\soc/cpu/pcpi_rs1 [5]),
    .Y(\soc/cpu/_02636_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07100_  (.A(\soc/cpu/decoded_imm[4] ),
    .B(\soc/cpu/pcpi_rs1 [4]),
    .Y(\soc/cpu/_02637_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07101_  (.A(\soc/cpu/decoded_imm[3] ),
    .B(\soc/cpu/pcpi_rs1 [3]),
    .Y(\soc/cpu/_02638_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07102_  (.A(\soc/cpu/decoded_imm[2] ),
    .B(\soc/cpu/pcpi_rs1 [2]),
    .X(\soc/cpu/_02639_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07103_  (.A(\soc/cpu/decoded_imm[2] ),
    .B(\soc/cpu/pcpi_rs1 [2]),
    .Y(\soc/cpu/_02640_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07104_  (.A(\soc/cpu/_02639_ ),
    .B(\soc/cpu/_02640_ ),
    .Y(\soc/cpu/_02641_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07105_  (.A(\soc/cpu/pcpi_rs1 [0]),
    .B(\soc/cpu/decoded_imm[0] ),
    .Y(\soc/cpu/_02642_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_07106_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/decoded_imm[1] ),
    .Y(\soc/cpu/_02643_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07107_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/decoded_imm[1] ),
    .Y(\soc/cpu/_02644_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07108_  (.A1(\soc/cpu/_02642_ ),
    .A2(\soc/cpu/_02643_ ),
    .B1(\soc/cpu/_02644_ ),
    .Y(\soc/cpu/_02645_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07109_  (.A(\soc/cpu/decoded_imm[3] ),
    .B(\soc/cpu/pcpi_rs1 [3]),
    .X(\soc/cpu/_02646_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_07110_  (.A1(\soc/cpu/_02641_ ),
    .A2(\soc/cpu/_02645_ ),
    .B1(\soc/cpu/_02646_ ),
    .C1(\soc/cpu/_02639_ ),
    .Y(\soc/cpu/_02647_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07111_  (.A(\soc/cpu/decoded_imm[4] ),
    .B(\soc/cpu/pcpi_rs1 [4]),
    .Y(\soc/cpu/_02648_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07112_  (.A(\soc/cpu/decoded_imm[5] ),
    .B(\soc/cpu/pcpi_rs1 [5]),
    .Y(\soc/cpu/_02649_ ));
 sky130_fd_sc_hd__o311a_1 \soc/cpu/_07113_  (.A1(\soc/cpu/_02637_ ),
    .A2(\soc/cpu/_02638_ ),
    .A3(\soc/cpu/_02647_ ),
    .B1(\soc/cpu/_02648_ ),
    .C1(\soc/cpu/_02649_ ),
    .X(\soc/cpu/_02650_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07114_  (.A(\soc/cpu/decoded_imm[6] ),
    .B(\soc/cpu/pcpi_rs1 [6]),
    .Y(\soc/cpu/_02651_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07115_  (.A(\soc/cpu/decoded_imm[7] ),
    .B(\soc/cpu/pcpi_rs1 [7]),
    .Y(\soc/cpu/_02652_ ));
 sky130_fd_sc_hd__o311a_1 \soc/cpu/_07116_  (.A1(\soc/cpu/_02635_ ),
    .A2(\soc/cpu/_02636_ ),
    .A3(\soc/cpu/_02650_ ),
    .B1(\soc/cpu/_02651_ ),
    .C1(\soc/cpu/_02652_ ),
    .X(\soc/cpu/_02653_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07117_  (.A(\soc/cpu/decoded_imm[8] ),
    .B(\soc/cpu/pcpi_rs1 [8]),
    .Y(\soc/cpu/_02654_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07118_  (.A(\soc/cpu/decoded_imm[9] ),
    .B(\soc/cpu/pcpi_rs1 [9]),
    .Y(\soc/cpu/_02655_ ));
 sky130_fd_sc_hd__o311ai_4 \soc/cpu/_07119_  (.A1(\soc/cpu/_02633_ ),
    .A2(\soc/cpu/_02634_ ),
    .A3(\soc/cpu/_02653_ ),
    .B1(\soc/cpu/_02654_ ),
    .C1(\soc/cpu/_02655_ ),
    .Y(\soc/cpu/_02656_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_07120_  (.A(\soc/cpu/decoded_imm[11] ),
    .B(\soc/cpu/pcpi_rs1 [11]),
    .X(\soc/cpu/_02657_ ));
 sky130_fd_sc_hd__a311oi_4 \soc/cpu/_07121_  (.A1(\soc/cpu/_02631_ ),
    .A2(\soc/cpu/_02632_ ),
    .A3(\soc/cpu/_02656_ ),
    .B1(\soc/cpu/_02629_ ),
    .C1(\soc/cpu/_02657_ ),
    .Y(\soc/cpu/_02658_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07122_  (.A(\soc/cpu/decoded_imm[12] ),
    .B(\soc/cpu/pcpi_rs1 [12]),
    .Y(\soc/cpu/_02659_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07123_  (.A(\soc/cpu/decoded_imm[13] ),
    .B(\soc/cpu/pcpi_rs1 [13]),
    .Y(\soc/cpu/_02660_ ));
 sky130_fd_sc_hd__o311ai_4 \soc/cpu/_07124_  (.A1(\soc/cpu/_02627_ ),
    .A2(\soc/cpu/_02628_ ),
    .A3(\soc/cpu/_02658_ ),
    .B1(\soc/cpu/_02659_ ),
    .C1(\soc/cpu/_02660_ ),
    .Y(\soc/cpu/_02661_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_07125_  (.A(\soc/cpu/decoded_imm[15] ),
    .B(\soc/cpu/pcpi_rs1 [15]),
    .X(\soc/cpu/_02662_ ));
 sky130_fd_sc_hd__a311oi_4 \soc/cpu/_07126_  (.A1(\soc/cpu/_02625_ ),
    .A2(\soc/cpu/_02626_ ),
    .A3(\soc/cpu/_02661_ ),
    .B1(\soc/cpu/_02623_ ),
    .C1(\soc/cpu/_02662_ ),
    .Y(\soc/cpu/_02663_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07127_  (.A(\soc/cpu/decoded_imm[16] ),
    .B(\soc/cpu/pcpi_rs1 [16]),
    .Y(\soc/cpu/_02664_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07128_  (.A(\soc/cpu/decoded_imm[17] ),
    .B(\soc/cpu/pcpi_rs1 [17]),
    .Y(\soc/cpu/_02665_ ));
 sky130_fd_sc_hd__o311ai_4 \soc/cpu/_07129_  (.A1(\soc/cpu/_02621_ ),
    .A2(\soc/cpu/_02622_ ),
    .A3(\soc/cpu/_02663_ ),
    .B1(\soc/cpu/_02664_ ),
    .C1(\soc/cpu/_02665_ ),
    .Y(\soc/cpu/_02666_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_07130_  (.A1(\soc/cpu/_02619_ ),
    .A2(\soc/cpu/_02620_ ),
    .A3(\soc/cpu/_02666_ ),
    .B1(\soc/cpu/_02617_ ),
    .Y(\soc/cpu/_02667_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07131_  (.A(\soc/cpu/decoded_imm[19] ),
    .B(\soc/cpu/pcpi_rs1 [19]),
    .Y(\soc/cpu/_02668_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07132_  (.A1(\soc/cpu/_02616_ ),
    .A2(\soc/cpu/_02667_ ),
    .B1(\soc/cpu/_02668_ ),
    .Y(\soc/cpu/_02669_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_07133_  (.A(\soc/cpu/decoded_imm[20] ),
    .B(\soc/cpu/pcpi_rs1 [20]),
    .C(\soc/cpu/_02669_ ),
    .X(\soc/cpu/_02670_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_07134_  (.A(\soc/cpu/decoded_imm[21] ),
    .B(\soc/cpu/pcpi_rs1 [21]),
    .C(\soc/cpu/_02670_ ),
    .X(\soc/cpu/_02671_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07135_  (.A(\soc/cpu/decoded_imm[22] ),
    .B(\soc/cpu/pcpi_rs1 [22]),
    .X(\soc/cpu/_02672_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_07136_  (.A1(\soc/cpu/_02615_ ),
    .A2(\soc/cpu/_02671_ ),
    .B1(\soc/cpu/_02672_ ),
    .Y(\soc/cpu/_02673_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07137_  (.A(\soc/cpu/decoded_imm[23] ),
    .B(\soc/cpu/pcpi_rs1 [23]),
    .Y(\soc/cpu/_02674_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07138_  (.A(\soc/cpu/decoded_imm[24] ),
    .B(\soc/cpu/pcpi_rs1 [24]),
    .Y(\soc/cpu/_02675_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07139_  (.A1(\soc/cpu/_02614_ ),
    .A2(\soc/cpu/_02673_ ),
    .B1(\soc/cpu/_02674_ ),
    .C1(\soc/cpu/_02675_ ),
    .Y(\soc/cpu/_02676_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_07140_  (.A1(\soc/cpu/decoded_imm[24] ),
    .A2(\soc/cpu/pcpi_rs1 [24]),
    .B1(\soc/cpu/_02676_ ),
    .Y(\soc/cpu/_02677_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07141_  (.A(\soc/cpu/decoded_imm[25] ),
    .B(\soc/cpu/pcpi_rs1 [25]),
    .Y(\soc/cpu/_02678_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07142_  (.A(\soc/cpu/decoded_imm[26] ),
    .B(\soc/cpu/pcpi_rs1 [26]),
    .Y(\soc/cpu/_02679_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07143_  (.A1(\soc/cpu/_02613_ ),
    .A2(\soc/cpu/_02677_ ),
    .B1(\soc/cpu/_02678_ ),
    .C1(\soc/cpu/_02679_ ),
    .Y(\soc/cpu/_02680_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07144_  (.A1(\soc/cpu/decoded_imm[26] ),
    .A2(\soc/cpu/pcpi_rs1 [26]),
    .B1(\soc/cpu/_02680_ ),
    .Y(\soc/cpu/_02681_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07145_  (.A(\soc/cpu/decoded_imm[27] ),
    .B(\soc/cpu/pcpi_rs1 [27]),
    .Y(\soc/cpu/_02682_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07146_  (.A1(\soc/cpu/_02612_ ),
    .A2(\soc/cpu/_02681_ ),
    .B1(\soc/cpu/_02682_ ),
    .Y(\soc/cpu/_02683_ ));
 sky130_fd_sc_hd__maj3_2 \soc/cpu/_07147_  (.A(\soc/cpu/decoded_imm[28] ),
    .B(\soc/cpu/pcpi_rs1 [28]),
    .C(\soc/cpu/_02683_ ),
    .X(\soc/cpu/_02684_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07148_  (.A(\soc/cpu/decoded_imm[29] ),
    .B(\soc/cpu/pcpi_rs1 [29]),
    .Y(\soc/cpu/_02685_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_07149_  (.A(\soc/cpu/_02685_ ),
    .Y(\soc/cpu/_02686_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07150_  (.A(\soc/cpu/decoded_imm[30] ),
    .B(\soc/cpu/pcpi_rs1 [30]),
    .X(\soc/cpu/_02687_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_07151_  (.A1(\soc/cpu/_02611_ ),
    .A2(\soc/cpu/_02684_ ),
    .B1(\soc/cpu/_02686_ ),
    .C1(\soc/cpu/_02687_ ),
    .Y(\soc/cpu/_02688_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07152_  (.A(\soc/cpu/decoded_imm[31] ),
    .B(\soc/cpu/pcpi_rs1 [31]),
    .Y(\soc/cpu/_02689_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_07153_  (.A1(\soc/cpu/_02610_ ),
    .A2(\soc/cpu/_02688_ ),
    .B1(\soc/cpu/_02689_ ),
    .X(\soc/cpu/_02690_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07154_  (.A1(\soc/cpu/_02610_ ),
    .A2(\soc/cpu/_02688_ ),
    .A3(\soc/cpu/_02689_ ),
    .B1(\soc/cpu/_00838_ ),
    .Y(\soc/cpu/_02691_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_07155_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/_01429_ ),
    .Y(\soc/cpu/_02692_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07157_  (.A(net343),
    .B(net353),
    .Y(\soc/cpu/_02694_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_07158_  (.A(\soc/cpu/cpuregs_raddr1[3] ),
    .B(net336),
    .C(net329),
    .Y(\soc/cpu/_02695_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_07159_  (.A(\soc/cpu/_02694_ ),
    .B(\soc/cpu/_02695_ ),
    .Y(\soc/cpu/_02696_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07161_  (.A(\soc/cpu/cpuregs_rdata1[31] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02698_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_16 \soc/cpu/_07162_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .SLEEP(\soc/cpu/instr_lui ),
    .X(\soc/cpu/_02699_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07164_  (.A(\soc/cpu/reg_pc[31] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_02701_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07165_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_02698_ ),
    .B1(\soc/cpu/_02701_ ),
    .Y(\soc/cpu/_02702_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07167_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/pcpi_rs1 [30]),
    .Y(\soc/cpu/_02704_ ));
 sky130_fd_sc_hd__nor4_4 \soc/cpu/_07168_  (.A(\soc/cpu/instr_sra ),
    .B(\soc/cpu/instr_srl ),
    .C(\soc/cpu/instr_srai ),
    .D(\soc/cpu/instr_srli ),
    .Y(\soc/cpu/_02705_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07170_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(\soc/cpu/_00936_ ),
    .B1(net155),
    .Y(\soc/cpu/_02707_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07171_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_02704_ ),
    .B1(\soc/cpu/_02707_ ),
    .Y(\soc/cpu/_02708_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07172_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_02702_ ),
    .B1(\soc/cpu/_02708_ ),
    .Y(\soc/cpu/_02709_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07173_  (.A(net47),
    .B(\soc/cpu/_02608_ ),
    .C(\soc/cpu/_02709_ ),
    .Y(\soc/cpu/_02710_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07174_  (.A1(\soc/cpu/_02690_ ),
    .A2(\soc/cpu/_02691_ ),
    .B1(\soc/cpu/_02710_ ),
    .Y(\soc/cpu/_02711_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07175_  (.A(\soc/cpu/_02609_ ),
    .B(\soc/cpu/_02711_ ),
    .Y(\soc/cpu/_00279_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07176_  (.A1(\soc/cpu/mem_la_read ),
    .A2(\soc/cpu/_00857_ ),
    .B1(\soc/cpu/_02352_ ),
    .Y(\soc/cpu/_02712_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07178_  (.A0(\soc/cpu/mem_la_addr [2]),
    .A1(\iomem_addr[2] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00503_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07179_  (.A0(\soc/cpu/mem_la_addr [3]),
    .A1(\iomem_addr[3] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00504_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07180_  (.A0(\soc/cpu/mem_la_addr [4]),
    .A1(\iomem_addr[4] ),
    .S(net51),
    .X(\soc/cpu/_00505_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07181_  (.A0(\soc/cpu/mem_la_addr [5]),
    .A1(\iomem_addr[5] ),
    .S(net51),
    .X(\soc/cpu/_00506_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07182_  (.A0(\soc/cpu/mem_la_addr [6]),
    .A1(\iomem_addr[6] ),
    .S(net51),
    .X(\soc/cpu/_00507_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07183_  (.A0(\soc/cpu/mem_la_addr [7]),
    .A1(\iomem_addr[7] ),
    .S(net51),
    .X(\soc/cpu/_00508_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07184_  (.A0(\soc/cpu/mem_la_addr [8]),
    .A1(\iomem_addr[8] ),
    .S(net51),
    .X(\soc/cpu/_00509_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07185_  (.A0(\soc/cpu/mem_la_addr [9]),
    .A1(\iomem_addr[9] ),
    .S(net51),
    .X(\soc/cpu/_00510_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07186_  (.A0(\soc/cpu/mem_la_addr [10]),
    .A1(\iomem_addr[10] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00511_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07187_  (.A0(\soc/cpu/mem_la_addr [11]),
    .A1(\iomem_addr[11] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00512_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07189_  (.A0(\soc/cpu/mem_la_addr [12]),
    .A1(\iomem_addr[12] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00513_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07190_  (.A0(\soc/cpu/mem_la_addr [13]),
    .A1(\iomem_addr[13] ),
    .S(net51),
    .X(\soc/cpu/_00514_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07191_  (.A0(\soc/cpu/mem_la_addr [14]),
    .A1(\iomem_addr[14] ),
    .S(net51),
    .X(\soc/cpu/_00515_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07192_  (.A0(\soc/cpu/mem_la_addr [15]),
    .A1(\iomem_addr[15] ),
    .S(net51),
    .X(\soc/cpu/_00516_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07193_  (.A0(\soc/cpu/mem_la_addr [16]),
    .A1(\iomem_addr[16] ),
    .S(net51),
    .X(\soc/cpu/_00517_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07194_  (.A0(\soc/cpu/mem_la_addr [17]),
    .A1(\iomem_addr[17] ),
    .S(net51),
    .X(\soc/cpu/_00518_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07195_  (.A0(\soc/cpu/mem_la_addr [18]),
    .A1(\iomem_addr[18] ),
    .S(net51),
    .X(\soc/cpu/_00519_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07196_  (.A0(\soc/cpu/mem_la_addr [19]),
    .A1(\iomem_addr[19] ),
    .S(net51),
    .X(\soc/cpu/_00520_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07197_  (.A0(\soc/cpu/mem_la_addr [20]),
    .A1(\iomem_addr[20] ),
    .S(net51),
    .X(\soc/cpu/_00521_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07198_  (.A0(\soc/cpu/mem_la_addr [21]),
    .A1(\iomem_addr[21] ),
    .S(net51),
    .X(\soc/cpu/_00522_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07200_  (.A0(\soc/cpu/mem_la_addr [22]),
    .A1(\iomem_addr[22] ),
    .S(net51),
    .X(\soc/cpu/_00523_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07201_  (.A0(\soc/cpu/mem_la_addr [23]),
    .A1(\iomem_addr[23] ),
    .S(net51),
    .X(\soc/cpu/_00524_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07202_  (.A0(\soc/cpu/mem_la_addr [24]),
    .A1(\iomem_addr[24] ),
    .S(net51),
    .X(\soc/cpu/_00525_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07203_  (.A0(\soc/cpu/mem_la_addr [25]),
    .A1(\iomem_addr[25] ),
    .S(net51),
    .X(\soc/cpu/_00526_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07204_  (.A0(\soc/cpu/mem_la_addr [26]),
    .A1(\iomem_addr[26] ),
    .S(net51),
    .X(\soc/cpu/_00527_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07205_  (.A0(\soc/cpu/mem_la_addr [27]),
    .A1(\iomem_addr[27] ),
    .S(net51),
    .X(\soc/cpu/_00528_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07206_  (.A0(\soc/cpu/mem_la_addr [28]),
    .A1(\iomem_addr[28] ),
    .S(net51),
    .X(\soc/cpu/_00529_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07207_  (.A0(\soc/cpu/mem_la_addr [29]),
    .A1(\iomem_addr[29] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00530_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07208_  (.A0(\soc/cpu/mem_la_addr [30]),
    .A1(\iomem_addr[30] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00531_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07209_  (.A0(\soc/cpu/mem_la_addr [31]),
    .A1(\iomem_addr[31] ),
    .S(\soc/cpu/_02712_ ),
    .X(\soc/cpu/_00532_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07210_  (.A(\soc/cpu/_01166_ ),
    .B(\soc/cpu/_01180_ ),
    .C(\soc/cpu/_02396_ ),
    .Y(\soc/cpu/_02716_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07211_  (.A1(\soc/cpu/_02387_ ),
    .A2(\soc/cpu/_02527_ ),
    .B1(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02717_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07212_  (.A(\soc/cpu/instr_lui ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02718_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07213_  (.A1(\soc/cpu/_02716_ ),
    .A2(\soc/cpu/_02717_ ),
    .B1(\soc/cpu/_02718_ ),
    .Y(\soc/cpu/_00533_ ));
 sky130_fd_sc_hd__a32o_1 \soc/cpu/_07214_  (.A1(\soc/cpu/_02412_ ),
    .A2(\soc/cpu/_02423_ ),
    .A3(\soc/cpu/_02424_ ),
    .B1(\soc/cpu/_02408_ ),
    .B2(\soc/cpu/instr_srai ),
    .X(\soc/cpu/_00534_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07215_  (.A(\soc/cpu/_01191_ ),
    .B(\soc/cpu/_01193_ ),
    .Y(\soc/cpu/_02719_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07216_  (.A(\soc/cpu/_01363_ ),
    .B(\soc/cpu/_01117_ ),
    .Y(\soc/cpu/_02720_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07217_  (.A(\soc/cpu/_01072_ ),
    .B(\soc/cpu/_01164_ ),
    .C(\soc/cpu/_01215_ ),
    .Y(\soc/cpu/_02721_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07218_  (.A(\soc/cpu/_01078_ ),
    .B(\soc/cpu/_02721_ ),
    .Y(\soc/cpu/_02722_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07219_  (.A1(\soc/cpu/_01124_ ),
    .A2(\soc/cpu/_02720_ ),
    .B1(\soc/cpu/_02722_ ),
    .Y(\soc/cpu/_02723_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07220_  (.A(\soc/cpu/_01233_ ),
    .B(\soc/cpu/_01211_ ),
    .Y(\soc/cpu/_02724_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07221_  (.A(\soc/cpu/_02529_ ),
    .B(\soc/cpu/_02724_ ),
    .Y(\soc/cpu/_02725_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07222_  (.A1(\soc/cpu/_01189_ ),
    .A2(\soc/cpu/_02723_ ),
    .B1(\soc/cpu/_02725_ ),
    .Y(\soc/cpu/_02726_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07223_  (.A1(\soc/cpu/_01215_ ),
    .A2(\soc/cpu/_01378_ ),
    .B1(\soc/cpu/_01081_ ),
    .Y(\soc/cpu/_02727_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07224_  (.A(\soc/cpu/_01233_ ),
    .B(\soc/cpu/_02727_ ),
    .Y(\soc/cpu/_02728_ ));
 sky130_fd_sc_hd__or4_2 \soc/cpu/_07225_  (.A(\soc/cpu/_01279_ ),
    .B(\soc/cpu/_02719_ ),
    .C(\soc/cpu/_02726_ ),
    .D(\soc/cpu/_02728_ ),
    .X(\soc/cpu/_02729_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07226_  (.A(\soc/cpu/_01212_ ),
    .B(\soc/cpu/_02729_ ),
    .Y(\soc/cpu/_02730_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07227_  (.A1(\soc/cpu/_01169_ ),
    .A2(\soc/cpu/_02441_ ),
    .B1(\soc/cpu/_02463_ ),
    .Y(\soc/cpu/_02731_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07228_  (.A1(\soc/cpu/cpuregs_raddr1[0] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02731_ ),
    .Y(\soc/cpu/_02732_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07229_  (.A1(\soc/cpu/_02446_ ),
    .A2(\soc/cpu/_02730_ ),
    .B1(\soc/cpu/_02732_ ),
    .Y(\soc/cpu/_00535_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07230_  (.A(\soc/cpu/_01169_ ),
    .B(\soc/cpu/_01155_ ),
    .Y(\soc/cpu/_02733_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07231_  (.A1(\soc/cpu/_01166_ ),
    .A2(\soc/cpu/_02398_ ),
    .B1(\soc/cpu/_02733_ ),
    .B2(\soc/cpu/_01192_ ),
    .C1(\soc/cpu/_02729_ ),
    .C2(\soc/cpu/_01137_ ),
    .Y(\soc/cpu/_02734_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_07232_  (.A1(\soc/cpu/_01237_ ),
    .A2(\soc/cpu/_02734_ ),
    .B1(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02735_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07233_  (.A1(\soc/cpu/_01342_ ),
    .A2(\soc/cpu/_02441_ ),
    .B1(\soc/cpu/_02463_ ),
    .Y(\soc/cpu/_02736_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/_07234_  (.A1(\soc/cpu/cpuregs_raddr1[1] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02735_ ),
    .C1(\soc/cpu/_02736_ ),
    .X(\soc/cpu/_00536_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07235_  (.A(\soc/cpu/_01140_ ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02737_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07236_  (.A1(\soc/cpu/cpuregs_raddr1[2] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02441_ ),
    .B2(\soc/cpu/_02480_ ),
    .C1(\soc/cpu/_02729_ ),
    .C2(\soc/cpu/_02737_ ),
    .Y(\soc/cpu/_02738_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_07237_  (.A(\soc/cpu/_02738_ ),
    .Y(\soc/cpu/_00537_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07238_  (.A(\soc/cpu/_00738_ ),
    .B(\soc/cpu/_01351_ ),
    .Y(\soc/cpu/_02739_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07239_  (.A1(\soc/cpu/_02441_ ),
    .A2(\soc/cpu/_02739_ ),
    .B1(\soc/cpu/_02726_ ),
    .B2(\soc/cpu/_01228_ ),
    .C1(\soc/cpu/_02719_ ),
    .Y(\soc/cpu/_02740_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07240_  (.A(\soc/cpu/_01279_ ),
    .B(\soc/cpu/_02446_ ),
    .C(\soc/cpu/_02728_ ),
    .Y(\soc/cpu/_02741_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07241_  (.A(\soc/cpu/cpuregs_raddr1[3] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02742_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07242_  (.A1(\soc/cpu/_02740_ ),
    .A2(\soc/cpu/_02741_ ),
    .B1(\soc/cpu/_02742_ ),
    .Y(\soc/cpu/_00538_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07243_  (.A(\soc/cpu/_00827_ ),
    .B(\soc/cpu/_01354_ ),
    .C(\soc/cpu/_02441_ ),
    .Y(\soc/cpu/_02743_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07244_  (.A1(\soc/cpu/_01118_ ),
    .A2(\soc/cpu/_01177_ ),
    .A3(\soc/cpu/_02404_ ),
    .B1(\soc/cpu/_01189_ ),
    .Y(\soc/cpu/_02744_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07245_  (.A1(\soc/cpu/_02724_ ),
    .A2(\soc/cpu/_02744_ ),
    .B1(\soc/cpu/_01130_ ),
    .Y(\soc/cpu/_02745_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07246_  (.A(\soc/cpu/cpuregs_raddr1[4] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02746_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07247_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02743_ ),
    .A3(\soc/cpu/_02745_ ),
    .B1(\soc/cpu/_02746_ ),
    .Y(\soc/cpu/_00539_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07248_  (.A1(\soc/cpu/_01080_ ),
    .A2(\soc/cpu/_02721_ ),
    .B1(\soc/cpu/_01189_ ),
    .Y(\soc/cpu/_02747_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07249_  (.A(\soc/cpu/_01081_ ),
    .B(\soc/cpu/_01215_ ),
    .C(\soc/cpu/_01166_ ),
    .Y(\soc/cpu/_02748_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_07250_  (.A1(\soc/cpu/_01193_ ),
    .A2(\soc/cpu/_01280_ ),
    .B1(\soc/cpu/_02748_ ),
    .B2(\soc/cpu/_01378_ ),
    .Y(\soc/cpu/_02749_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07251_  (.A1(\soc/cpu/_02747_ ),
    .A2(\soc/cpu/_02749_ ),
    .B1(\soc/cpu/_01110_ ),
    .Y(\soc/cpu/_02750_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07252_  (.A(\soc/cpu/cpuregs_raddr2[0] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02751_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07253_  (.A1(\soc/cpu/_02470_ ),
    .A2(\soc/cpu/_02750_ ),
    .B1(\soc/cpu/_02751_ ),
    .Y(\soc/cpu/_00540_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_07254_  (.A(\soc/cpu/cpuregs_raddr2[1] ),
    .Y(\soc/cpu/_02752_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_07255_  (.A1(\soc/cpu/_02747_ ),
    .A2(\soc/cpu/_02749_ ),
    .B1(\soc/cpu/_01116_ ),
    .C1(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02753_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_07256_  (.A1(\soc/cpu/_02752_ ),
    .A2(\soc/cpu/_01588_ ),
    .B1(\soc/cpu/_02449_ ),
    .C1(\soc/cpu/_02753_ ),
    .Y(\soc/cpu/_00541_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_07257_  (.A1(\soc/cpu/_01117_ ),
    .A2(\soc/cpu/_02404_ ),
    .B1(\soc/cpu/_01080_ ),
    .X(\soc/cpu/_02754_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07258_  (.A(\soc/cpu/_01189_ ),
    .B(\soc/cpu/_02754_ ),
    .Y(\soc/cpu/_02755_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07259_  (.A1(\soc/cpu/_02749_ ),
    .A2(\soc/cpu/_02755_ ),
    .B1(\soc/cpu/_02452_ ),
    .Y(\soc/cpu/_02756_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_07260_  (.A1(\soc/cpu/_01411_ ),
    .A2(\soc/cpu/_01588_ ),
    .B1(\soc/cpu/_02450_ ),
    .C1(\soc/cpu/_02756_ ),
    .Y(\soc/cpu/_00542_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07261_  (.A(\soc/cpu/_01130_ ),
    .B(\soc/cpu/_02748_ ),
    .Y(\soc/cpu/_02757_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07262_  (.A1(\soc/cpu/_02755_ ),
    .A2(\soc/cpu/_02757_ ),
    .B1(\soc/cpu/_01210_ ),
    .Y(\soc/cpu/_02758_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_07263_  (.A(\soc/cpu/_01290_ ),
    .B(\soc/cpu/_02446_ ),
    .C(\soc/cpu/_02388_ ),
    .D(\soc/cpu/_02456_ ),
    .Y(\soc/cpu/_02759_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07264_  (.A(\soc/cpu/cpuregs_raddr2[3] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02760_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07265_  (.A1(\soc/cpu/_02758_ ),
    .A2(\soc/cpu/_02759_ ),
    .B1(\soc/cpu/_02760_ ),
    .Y(\soc/cpu/_00543_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07266_  (.A1(\soc/cpu/_02747_ ),
    .A2(\soc/cpu/_02757_ ),
    .B1(\soc/cpu/_01289_ ),
    .Y(\soc/cpu/_02761_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07267_  (.A(\soc/cpu/cpuregs_raddr2[4] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02762_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07268_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02458_ ),
    .A3(\soc/cpu/_02761_ ),
    .B1(\soc/cpu/_02762_ ),
    .Y(\soc/cpu/_00544_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07269_  (.A(\soc/cpu/is_sb_sh_sw ),
    .B(\soc/cpu/mem_rdata_q[7] ),
    .C(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02763_ ));
 sky130_fd_sc_hd__or3_2 \soc/cpu/_07270_  (.A(\soc/cpu/instr_jalr ),
    .B(\soc/cpu/is_lb_lh_lw_lbu_lhu ),
    .C(net697),
    .X(\soc/cpu/_02764_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07272_  (.A(\soc/cpu/mem_rdata_q[20] ),
    .B(\soc/cpu/_02411_ ),
    .C(\soc/cpu/_02764_ ),
    .Y(\soc/cpu/_02766_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07274_  (.A(\soc/cpu/decoded_imm[0] ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02768_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07275_  (.A(\soc/cpu/_02763_ ),
    .B(\soc/cpu/_02766_ ),
    .C(\soc/cpu/_02768_ ),
    .Y(\soc/cpu/_00545_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_07278_  (.A(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .B(\soc/cpu/is_sb_sh_sw ),
    .X(\soc/cpu/_02771_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07279_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[1] ),
    .B1(\soc/cpu/_02771_ ),
    .B2(\soc/cpu/mem_rdata_q[8] ),
    .C1(\soc/cpu/_02764_ ),
    .C2(\soc/cpu/mem_rdata_q[21] ),
    .Y(\soc/cpu/_02772_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07280_  (.A(\soc/cpu/decoded_imm[1] ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02773_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07281_  (.A1(\soc/cpu/_02408_ ),
    .A2(\soc/cpu/_02772_ ),
    .B1(\soc/cpu/_02773_ ),
    .Y(\soc/cpu/_00546_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07282_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[2] ),
    .B1(\soc/cpu/_02771_ ),
    .B2(\soc/cpu/mem_rdata_q[9] ),
    .C1(\soc/cpu/_02764_ ),
    .C2(\soc/cpu/mem_rdata_q[22] ),
    .Y(\soc/cpu/_02774_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07283_  (.A(\soc/cpu/decoded_imm[2] ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02775_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07284_  (.A1(\soc/cpu/_02408_ ),
    .A2(\soc/cpu/_02774_ ),
    .B1(\soc/cpu/_02775_ ),
    .Y(\soc/cpu/_00547_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07285_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[3] ),
    .B1(\soc/cpu/_02764_ ),
    .B2(\soc/cpu/mem_rdata_q[23] ),
    .C1(\soc/cpu/_02771_ ),
    .C2(\soc/cpu/mem_rdata_q[10] ),
    .Y(\soc/cpu/_02776_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07286_  (.A(\soc/cpu/decoded_imm[3] ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02777_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07287_  (.A1(\soc/cpu/_02408_ ),
    .A2(\soc/cpu/_02776_ ),
    .B1(\soc/cpu/_02777_ ),
    .Y(\soc/cpu/_00548_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07288_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[4] ),
    .B1(\soc/cpu/_02764_ ),
    .B2(\soc/cpu/mem_rdata_q[24] ),
    .C1(\soc/cpu/_02771_ ),
    .C2(\soc/cpu/mem_rdata_q[11] ),
    .Y(\soc/cpu/_02778_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07289_  (.A(\soc/cpu/decoded_imm[4] ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02779_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07290_  (.A1(\soc/cpu/_02408_ ),
    .A2(\soc/cpu/_02778_ ),
    .B1(\soc/cpu/_02779_ ),
    .Y(\soc/cpu/_00549_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_07291_  (.A(\soc/cpu/_02764_ ),
    .B(\soc/cpu/_02771_ ),
    .X(\soc/cpu/_02780_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07293_  (.A(\soc/cpu/mem_rdata_q[25] ),
    .B(\soc/cpu/_02411_ ),
    .C(\soc/cpu/_02780_ ),
    .Y(\soc/cpu/_02782_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07294_  (.A(\soc/cpu/decoded_imm[5] ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02783_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07295_  (.A(\soc/cpu/instr_jal ),
    .B(\soc/cpu/decoded_imm_j[5] ),
    .C(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02784_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07296_  (.A(\soc/cpu/_02782_ ),
    .B(\soc/cpu/_02783_ ),
    .C(\soc/cpu/_02784_ ),
    .Y(\soc/cpu/_00550_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07297_  (.A(\soc/cpu/decoded_imm[6] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02785_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07298_  (.A1(\soc/cpu/instr_jal ),
    .A2(net964),
    .B1(\soc/cpu/_02780_ ),
    .B2(\soc/cpu/mem_rdata_q[26] ),
    .C1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02786_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07299_  (.A(\soc/cpu/_02785_ ),
    .B(net965),
    .Y(\soc/cpu/_00551_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07300_  (.A(\soc/cpu/decoded_imm[7] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02787_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07301_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[7] ),
    .B1(\soc/cpu/_02780_ ),
    .B2(\soc/cpu/mem_rdata_q[27] ),
    .C1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02788_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07302_  (.A(\soc/cpu/_02787_ ),
    .B(\soc/cpu/_02788_ ),
    .Y(\soc/cpu/_00552_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07303_  (.A(\soc/cpu/decoded_imm[8] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02789_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07304_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[8] ),
    .B1(\soc/cpu/_02780_ ),
    .B2(\soc/cpu/mem_rdata_q[28] ),
    .C1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02790_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07305_  (.A(\soc/cpu/_02789_ ),
    .B(\soc/cpu/_02790_ ),
    .Y(\soc/cpu/_00553_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07306_  (.A(\soc/cpu/decoded_imm[9] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02791_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07307_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[9] ),
    .B1(\soc/cpu/_02780_ ),
    .B2(\soc/cpu/mem_rdata_q[29] ),
    .C1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02792_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07308_  (.A(\soc/cpu/_02791_ ),
    .B(\soc/cpu/_02792_ ),
    .Y(\soc/cpu/_00554_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07309_  (.A(\soc/cpu/decoded_imm[10] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02793_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_07310_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[10] ),
    .B1(\soc/cpu/_02780_ ),
    .B2(\soc/cpu/mem_rdata_q[30] ),
    .C1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02794_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07311_  (.A(\soc/cpu/_02793_ ),
    .B(\soc/cpu/_02794_ ),
    .Y(\soc/cpu/_00555_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07312_  (.A1(\soc/cpu/mem_rdata_q[31] ),
    .A2(\soc/cpu/_02764_ ),
    .B1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02795_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_07313_  (.A1(\soc/cpu/is_sb_sh_sw ),
    .A2(\soc/cpu/mem_rdata_q[31] ),
    .B1(\soc/cpu/mem_rdata_q[7] ),
    .B2(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .C1(\soc/cpu/instr_jal ),
    .C2(\soc/cpu/decoded_imm_j[11] ),
    .Y(\soc/cpu/_02796_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07315_  (.A(\soc/cpu/decoded_imm[11] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02798_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07316_  (.A1(\soc/cpu/_02795_ ),
    .A2(\soc/cpu/_02796_ ),
    .B1(\soc/cpu/_02798_ ),
    .Y(\soc/cpu/_00556_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_07317_  (.A1(\soc/cpu/mem_rdata_q[31] ),
    .A2(\soc/cpu/_02780_ ),
    .B1(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02799_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07319_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[12] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(\soc/cpu/mem_rdata_q[12] ),
    .Y(\soc/cpu/_02801_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07320_  (.A(\soc/cpu/decoded_imm[12] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02802_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07321_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02801_ ),
    .B1(\soc/cpu/_02802_ ),
    .Y(\soc/cpu/_00557_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07322_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[13] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(net956),
    .Y(\soc/cpu/_02803_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07323_  (.A(\soc/cpu/decoded_imm[13] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02804_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07324_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02803_ ),
    .B1(\soc/cpu/_02804_ ),
    .Y(\soc/cpu/_00558_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07325_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[14] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(net852),
    .Y(\soc/cpu/_02805_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07326_  (.A(\soc/cpu/decoded_imm[14] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02806_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07327_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02805_ ),
    .B1(\soc/cpu/_02806_ ),
    .Y(\soc/cpu/_00559_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07328_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[15] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(\soc/cpu/mem_rdata_q[15] ),
    .Y(\soc/cpu/_02807_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07329_  (.A(\soc/cpu/decoded_imm[15] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02808_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07330_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02807_ ),
    .B1(\soc/cpu/_02808_ ),
    .Y(\soc/cpu/_00560_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07331_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[16] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(\soc/cpu/mem_rdata_q[16] ),
    .Y(\soc/cpu/_02809_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07332_  (.A(\soc/cpu/decoded_imm[16] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02810_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07333_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02809_ ),
    .B1(\soc/cpu/_02810_ ),
    .Y(\soc/cpu/_00561_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07334_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[17] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(\soc/cpu/mem_rdata_q[17] ),
    .Y(\soc/cpu/_02811_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07335_  (.A(\soc/cpu/decoded_imm[17] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02812_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07336_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02811_ ),
    .B1(\soc/cpu/_02812_ ),
    .Y(\soc/cpu/_00562_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07337_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[18] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(\soc/cpu/mem_rdata_q[18] ),
    .Y(\soc/cpu/_02813_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07339_  (.A(\soc/cpu/decoded_imm[18] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02815_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07340_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02813_ ),
    .B1(\soc/cpu/_02815_ ),
    .Y(\soc/cpu/_00563_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_07341_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[19] ),
    .B1(\soc/cpu/_00878_ ),
    .B2(\soc/cpu/mem_rdata_q[19] ),
    .Y(\soc/cpu/_02816_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07342_  (.A(\soc/cpu/decoded_imm[19] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02817_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07343_  (.A1(\soc/cpu/_02799_ ),
    .A2(\soc/cpu/_02816_ ),
    .B1(\soc/cpu/_02817_ ),
    .Y(\soc/cpu/_00564_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07345_  (.A(\soc/cpu/mem_rdata_q[20] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02819_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_07348_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[20] ),
    .B1_N(\soc/cpu/_02799_ ),
    .Y(\soc/cpu/_02822_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07349_  (.A(\soc/cpu/decoded_imm[20] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02823_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07350_  (.A1(\soc/cpu/_02819_ ),
    .A2(\soc/cpu/_02822_ ),
    .B1(\soc/cpu/_02823_ ),
    .Y(\soc/cpu/_00565_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07352_  (.A(\soc/cpu/mem_rdata_q[21] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02825_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07353_  (.A(\soc/cpu/decoded_imm[21] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02826_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07354_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02825_ ),
    .B1(\soc/cpu/_02826_ ),
    .Y(\soc/cpu/_00566_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07355_  (.A(\soc/cpu/mem_rdata_q[22] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02827_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07356_  (.A(\soc/cpu/decoded_imm[22] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02828_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07357_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02827_ ),
    .B1(\soc/cpu/_02828_ ),
    .Y(\soc/cpu/_00567_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07358_  (.A(\soc/cpu/mem_rdata_q[23] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02829_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07359_  (.A(\soc/cpu/decoded_imm[23] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02830_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07360_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02829_ ),
    .B1(\soc/cpu/_02830_ ),
    .Y(\soc/cpu/_00568_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07361_  (.A(net957),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02831_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07362_  (.A(\soc/cpu/decoded_imm[24] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02832_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07363_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02831_ ),
    .B1(\soc/cpu/_02832_ ),
    .Y(\soc/cpu/_00569_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07364_  (.A(\soc/cpu/mem_rdata_q[25] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02833_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07365_  (.A(\soc/cpu/decoded_imm[25] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02834_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07366_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02833_ ),
    .B1(\soc/cpu/_02834_ ),
    .Y(\soc/cpu/_00570_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07367_  (.A(\soc/cpu/mem_rdata_q[26] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02835_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07368_  (.A(\soc/cpu/decoded_imm[26] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02836_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07369_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02835_ ),
    .B1(\soc/cpu/_02836_ ),
    .Y(\soc/cpu/_00571_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07370_  (.A(net875),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02837_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07371_  (.A(\soc/cpu/decoded_imm[27] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02838_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07372_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02837_ ),
    .B1(\soc/cpu/_02838_ ),
    .Y(\soc/cpu/_00572_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07373_  (.A(\soc/cpu/mem_rdata_q[28] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02839_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07374_  (.A(\soc/cpu/decoded_imm[28] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02840_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07375_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02839_ ),
    .B1(\soc/cpu/_02840_ ),
    .Y(\soc/cpu/_00573_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07376_  (.A(\soc/cpu/mem_rdata_q[29] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02841_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07377_  (.A(\soc/cpu/decoded_imm[29] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02842_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07378_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02841_ ),
    .B1(\soc/cpu/_02842_ ),
    .Y(\soc/cpu/_00574_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07379_  (.A(\soc/cpu/mem_rdata_q[30] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02843_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07380_  (.A(\soc/cpu/decoded_imm[30] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02844_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07381_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02843_ ),
    .B1(\soc/cpu/_02844_ ),
    .Y(\soc/cpu/_00575_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07382_  (.A(\soc/cpu/mem_rdata_q[31] ),
    .B(\soc/cpu/_00878_ ),
    .Y(\soc/cpu/_02845_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07383_  (.A(\soc/cpu/decoded_imm[31] ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_02846_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07384_  (.A1(\soc/cpu/_02822_ ),
    .A2(\soc/cpu/_02845_ ),
    .B1(\soc/cpu/_02846_ ),
    .Y(\soc/cpu/_00576_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07385_  (.A1(net697),
    .A2(\soc/cpu/_02508_ ),
    .B1(\soc/cpu/instr_jalr ),
    .Y(\soc/cpu/_02847_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07386_  (.A(\soc/cpu/is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02848_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07387_  (.A1(\soc/cpu/_02408_ ),
    .A2(net698),
    .B1(\soc/cpu/_02848_ ),
    .Y(\soc/cpu/_00577_ ));
 sky130_fd_sc_hd__a41oi_2 \soc/cpu/_07388_  (.A1(\soc/cpu/_01210_ ),
    .A2(\soc/cpu/_01095_ ),
    .A3(\soc/cpu/_01102_ ),
    .A4(\soc/cpu/_02386_ ),
    .B1(\soc/cpu/_01281_ ),
    .Y(\soc/cpu/_02849_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07389_  (.A(\soc/cpu/is_sb_sh_sw ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02850_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07390_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02849_ ),
    .B1(\soc/cpu/_02850_ ),
    .Y(\soc/cpu/_00578_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07391_  (.A(\soc/cpu/compressed_instr ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02851_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07392_  (.A(\soc/cpu/_02448_ ),
    .B(\soc/cpu/_02851_ ),
    .Y(\soc/cpu/_00580_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07393_  (.A(\soc/cpu/instr_lb ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02852_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07394_  (.A1(\soc/cpu/_02516_ ),
    .A2(\soc/cpu/_02519_ ),
    .B1(\soc/cpu/_02852_ ),
    .Y(\soc/cpu/_00619_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07395_  (.A(\soc/cpu/instr_lw ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02853_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07396_  (.A1(\soc/cpu/_02491_ ),
    .A2(\soc/cpu/_02519_ ),
    .B1(\soc/cpu/_02853_ ),
    .Y(\soc/cpu/_00620_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07398_  (.A(\soc/cpu/instr_rdinstr ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02855_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07399_  (.A1(\soc/cpu/_02498_ ),
    .A2(\soc/cpu/_02504_ ),
    .B1(\soc/cpu/_02855_ ),
    .Y(\soc/cpu/_00623_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07400_  (.A(\soc/cpu/_01205_ ),
    .B(\soc/cpu/_01224_ ),
    .Y(\soc/cpu/_02856_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_07401_  (.A(\soc/cpu/_02446_ ),
    .B(\soc/cpu/_02437_ ),
    .C(\soc/cpu/_02440_ ),
    .D(\soc/cpu/_02856_ ),
    .Y(\soc/cpu/_02857_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_07402_  (.A1(\soc/cpu/instr_waitirq ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02857_ ),
    .X(\soc/cpu/_00624_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07404_  (.A(\soc/cpu/instr_timer ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02859_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07405_  (.A(\soc/cpu/_02418_ ),
    .B(\soc/cpu/_02431_ ),
    .C(\soc/cpu/_02486_ ),
    .Y(\soc/cpu/_02860_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07406_  (.A(\soc/cpu/_02859_ ),
    .B(\soc/cpu/_02860_ ),
    .Y(\soc/cpu/_00625_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07407_  (.A1(\soc/cpu/_01235_ ),
    .A2(\soc/cpu/_02397_ ),
    .B1(\soc/cpu/_01233_ ),
    .Y(\soc/cpu/_02861_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07408_  (.A(\soc/cpu/_01358_ ),
    .B(\soc/cpu/_02720_ ),
    .C(\soc/cpu/_02722_ ),
    .Y(\soc/cpu/_02862_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07409_  (.A1(\soc/cpu/_00826_ ),
    .A2(\soc/cpu/_02862_ ),
    .B1(\soc/cpu/_00738_ ),
    .Y(\soc/cpu/_02863_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07410_  (.A(\soc/cpu/_02861_ ),
    .B(\soc/cpu/_02863_ ),
    .Y(\soc/cpu/_02864_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07411_  (.A1(\soc/cpu/_01233_ ),
    .A2(\soc/cpu/_02727_ ),
    .B1(\soc/cpu/_02864_ ),
    .Y(\soc/cpu/_02865_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_07412_  (.A1(\soc/cpu/_01193_ ),
    .A2(\soc/cpu/_01208_ ),
    .B1(\soc/cpu/_01248_ ),
    .B2(\soc/cpu/_01078_ ),
    .Y(\soc/cpu/_02866_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07413_  (.A1(\soc/cpu/_01124_ ),
    .A2(\soc/cpu/_02529_ ),
    .B1(\soc/cpu/_02865_ ),
    .B2(\soc/cpu/_01212_ ),
    .C1(\soc/cpu/_02866_ ),
    .Y(\soc/cpu/_02867_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07414_  (.A(\soc/cpu/decoded_rd[0] ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02868_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07415_  (.A1(\soc/cpu/_02446_ ),
    .A2(\soc/cpu/_02867_ ),
    .B1(\soc/cpu/_02868_ ),
    .Y(\soc/cpu/_00626_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07416_  (.A(\soc/cpu/decoded_rd[1] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02869_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07417_  (.A1(\soc/cpu/_01198_ ),
    .A2(\soc/cpu/_01242_ ),
    .B1(\soc/cpu/_02865_ ),
    .B2(\soc/cpu/_01137_ ),
    .C1(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02870_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07418_  (.A(\soc/cpu/_02869_ ),
    .B(\soc/cpu/_02870_ ),
    .Y(\soc/cpu/_00627_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07419_  (.A(\soc/cpu/_01102_ ),
    .B(\soc/cpu/_01404_ ),
    .C(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02871_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_07420_  (.A1(\soc/cpu/decoded_rd[2] ),
    .A2(\soc/cpu/_02446_ ),
    .B1(\soc/cpu/_02737_ ),
    .B2(\soc/cpu/_02865_ ),
    .C1(\soc/cpu/_02871_ ),
    .X(\soc/cpu/_00628_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07421_  (.A(\soc/cpu/_01152_ ),
    .B(\soc/cpu/_02727_ ),
    .Y(\soc/cpu/_02872_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07422_  (.A1(\soc/cpu/_02728_ ),
    .A2(\soc/cpu/_02861_ ),
    .B1(\soc/cpu/_02872_ ),
    .Y(\soc/cpu/_02873_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07423_  (.A1(\soc/cpu/_01228_ ),
    .A2(\soc/cpu/_02863_ ),
    .B1(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02874_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07424_  (.A(\soc/cpu/decoded_rd[3] ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02875_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07425_  (.A1(\soc/cpu/_01404_ ),
    .A2(\soc/cpu/_02873_ ),
    .A3(\soc/cpu/_02874_ ),
    .B1(\soc/cpu/_02875_ ),
    .Y(\soc/cpu/_00629_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07426_  (.A(\soc/cpu/decoded_rd[4] ),
    .B(\soc/cpu/_02446_ ),
    .Y(\soc/cpu/_02876_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07427_  (.A1(\soc/cpu/_01171_ ),
    .A2(\soc/cpu/_02446_ ),
    .A3(\soc/cpu/_02864_ ),
    .B1(\soc/cpu/_02876_ ),
    .Y(\soc/cpu/_00630_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07428_  (.A(\soc/cpu/_01235_ ),
    .B(\soc/cpu/_01193_ ),
    .Y(\soc/cpu/_02877_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07429_  (.A(\soc/cpu/_01189_ ),
    .B(\soc/cpu/_01155_ ),
    .C(\soc/cpu/_01391_ ),
    .Y(\soc/cpu/_02878_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_07430_  (.A1(\soc/cpu/_00827_ ),
    .A2(\soc/cpu/_01117_ ),
    .B1(\soc/cpu/_02877_ ),
    .B2(\soc/cpu/_01064_ ),
    .C1(\soc/cpu/_02878_ ),
    .Y(\soc/cpu/_02879_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07431_  (.A(\soc/cpu/is_lb_lh_lw_lbu_lhu ),
    .B(\soc/cpu/_01588_ ),
    .Y(\soc/cpu/_02880_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07432_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_02879_ ),
    .B1(\soc/cpu/_02880_ ),
    .Y(\soc/cpu/_00631_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07433_  (.A(\soc/cpu/is_sll_srl_sra ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_02881_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07434_  (.A(net850),
    .B(\soc/cpu/_02411_ ),
    .C(\soc/cpu/_02426_ ),
    .Y(\soc/cpu/_02882_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07435_  (.A(\soc/cpu/_02881_ ),
    .B(\soc/cpu/_02882_ ),
    .Y(\soc/cpu/_00632_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07436_  (.A0(\soc/cpu/mem_la_wdata [0]),
    .A1(\iomem_wdata[0] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00633_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07438_  (.A(\iomem_wdata[1] ),
    .B(\soc/cpu/_02382_ ),
    .Y(\soc/cpu/_02884_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07439_  (.A1(\soc/cpu/_01521_ ),
    .A2(\soc/cpu/_02382_ ),
    .B1(\soc/cpu/_02884_ ),
    .Y(\soc/cpu/_00634_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07440_  (.A(net276),
    .B(\soc/cpu/_02382_ ),
    .Y(\soc/cpu/_02885_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07441_  (.A1(\soc/cpu/_01520_ ),
    .A2(\soc/cpu/_02382_ ),
    .B1(\soc/cpu/_02885_ ),
    .Y(\soc/cpu/_00635_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07442_  (.A(net268),
    .B(\soc/cpu/_02382_ ),
    .Y(\soc/cpu/_02886_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07443_  (.A1(\soc/cpu/_01519_ ),
    .A2(\soc/cpu/_02382_ ),
    .B1(\soc/cpu/_02886_ ),
    .Y(\soc/cpu/_00636_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07444_  (.A(\iomem_wdata[4] ),
    .B(\soc/cpu/_02382_ ),
    .Y(\soc/cpu/_02887_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07445_  (.A1(\soc/cpu/_01518_ ),
    .A2(\soc/cpu/_02382_ ),
    .B1(\soc/cpu/_02887_ ),
    .Y(\soc/cpu/_00637_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07446_  (.A(\iomem_wdata[5] ),
    .B(\soc/cpu/_02382_ ),
    .Y(\soc/cpu/_02888_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07447_  (.A1(\soc/cpu/_01517_ ),
    .A2(\soc/cpu/_02382_ ),
    .B1(\soc/cpu/_02888_ ),
    .Y(\soc/cpu/_00638_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07448_  (.A0(net776),
    .A1(\iomem_wdata[6] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00639_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07449_  (.A(\iomem_wdata[7] ),
    .B(\soc/cpu/_02382_ ),
    .Y(\soc/cpu/_02889_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07450_  (.A1(\soc/cpu/_01516_ ),
    .A2(\soc/cpu/_02382_ ),
    .B1(\soc/cpu/_02889_ ),
    .Y(\soc/cpu/_00640_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07451_  (.A0(\soc/cpu/mem_la_wdata [8]),
    .A1(\iomem_wdata[8] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00641_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07452_  (.A0(\soc/cpu/mem_la_wdata [9]),
    .A1(\iomem_wdata[9] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00642_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07453_  (.A0(\soc/cpu/mem_la_wdata [10]),
    .A1(\iomem_wdata[10] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00643_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07454_  (.A0(\soc/cpu/mem_la_wdata [11]),
    .A1(\iomem_wdata[11] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00644_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07456_  (.A0(\soc/cpu/mem_la_wdata [12]),
    .A1(\iomem_wdata[12] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00645_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07457_  (.A0(\soc/cpu/mem_la_wdata [13]),
    .A1(\iomem_wdata[13] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00646_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07458_  (.A0(\soc/cpu/mem_la_wdata [14]),
    .A1(\iomem_wdata[14] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00647_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07459_  (.A0(\soc/cpu/mem_la_wdata [15]),
    .A1(\iomem_wdata[15] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00648_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07460_  (.A0(\soc/cpu/mem_la_wdata [16]),
    .A1(\iomem_wdata[16] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00649_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07461_  (.A0(\soc/cpu/mem_la_wdata [17]),
    .A1(\iomem_wdata[17] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00650_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07462_  (.A0(\soc/cpu/mem_la_wdata [18]),
    .A1(\iomem_wdata[18] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00651_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07463_  (.A0(\soc/cpu/mem_la_wdata [19]),
    .A1(\iomem_wdata[19] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00652_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07464_  (.A0(\soc/cpu/mem_la_wdata [20]),
    .A1(\iomem_wdata[20] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00653_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07465_  (.A0(\soc/cpu/mem_la_wdata [21]),
    .A1(\iomem_wdata[21] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00654_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07467_  (.A0(\soc/cpu/mem_la_wdata [22]),
    .A1(\iomem_wdata[22] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00655_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07468_  (.A0(\soc/cpu/mem_la_wdata [23]),
    .A1(\iomem_wdata[23] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00656_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07469_  (.A0(\soc/cpu/mem_la_wdata [24]),
    .A1(\iomem_wdata[24] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00657_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07470_  (.A0(\soc/cpu/mem_la_wdata [25]),
    .A1(\iomem_wdata[25] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00658_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07471_  (.A0(\soc/cpu/mem_la_wdata [26]),
    .A1(\iomem_wdata[26] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00659_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07472_  (.A0(\soc/cpu/mem_la_wdata [27]),
    .A1(\iomem_wdata[27] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00660_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07473_  (.A0(\soc/cpu/mem_la_wdata [28]),
    .A1(\iomem_wdata[28] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00661_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07474_  (.A0(\soc/cpu/mem_la_wdata [29]),
    .A1(\iomem_wdata[29] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00662_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07475_  (.A0(\soc/cpu/mem_la_wdata [30]),
    .A1(\iomem_wdata[30] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00663_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_07476_  (.A0(\soc/cpu/mem_la_wdata [31]),
    .A1(\iomem_wdata[31] ),
    .S(\soc/cpu/_02382_ ),
    .X(\soc/cpu/_00664_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_07477_  (.A(\soc/cpu/_00744_ ),
    .B(\soc/cpu/_02351_ ),
    .C(\soc/cpu/_02352_ ),
    .X(\soc/cpu/_02892_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07478_  (.A1(\soc/cpu/mem_do_rinst ),
    .A2(\soc/cpu/_02367_ ),
    .A3(\soc/cpu/_02362_ ),
    .B1(\soc/cpu/_02369_ ),
    .Y(\soc/cpu/_02893_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07479_  (.A(\soc/cpu/_02364_ ),
    .B(\soc/cpu/_02366_ ),
    .C(\soc/cpu/_02892_ ),
    .D(\soc/cpu/_02893_ ),
    .Y(\soc/cpu/_02894_ ));
 sky130_fd_sc_hd__or4_1 \soc/cpu/_07480_  (.A(\soc/cpu/mem_do_rinst ),
    .B(\soc/cpu/mem_do_rdata ),
    .C(\soc/cpu/_02350_ ),
    .D(\soc/cpu/_02362_ ),
    .X(\soc/cpu/_02895_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07481_  (.A(\soc/cpu/mem_state[0] ),
    .B(\soc/cpu/_02894_ ),
    .Y(\soc/cpu/_02896_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07482_  (.A1(\soc/cpu/_02365_ ),
    .A2(\soc/cpu/_02894_ ),
    .A3(\soc/cpu/_02895_ ),
    .B1(\soc/cpu/_02896_ ),
    .Y(\soc/cpu/_00666_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07483_  (.A(\soc/cpu/mem_state[1] ),
    .B(\soc/cpu/_02894_ ),
    .Y(\soc/cpu/_02897_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07484_  (.A1(\soc/cpu/_02382_ ),
    .A2(\soc/cpu/_02894_ ),
    .A3(\soc/cpu/_02895_ ),
    .B1(\soc/cpu/_02897_ ),
    .Y(\soc/cpu/_00667_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07485_  (.A1(\soc/cpu/cpuregs_rdata2[0] ),
    .A2(\soc/cpu/_01414_ ),
    .B1(\soc/cpu/is_slli_srli_srai ),
    .Y(\soc/cpu/_02898_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_07486_  (.A(\soc/cpu/is_slli_srli_srai ),
    .SLEEP(\soc/cpu/cpuregs_raddr2[0] ),
    .X(\soc/cpu/_02899_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07488_  (.A(\soc/cpu/reg_sh[0] ),
    .B(\soc/cpu/_00937_ ),
    .Y(\soc/cpu/_02901_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07489_  (.A1(\soc/cpu/reg_sh[0] ),
    .A2(\soc/cpu/_01421_ ),
    .B1(\soc/cpu/_02901_ ),
    .Y(\soc/cpu/_02902_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07490_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/_02898_ ),
    .A3(\soc/cpu/_02899_ ),
    .B1(\soc/cpu/_02902_ ),
    .Y(\soc/cpu/_00668_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07491_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/reg_sh[1] ),
    .C(\soc/cpu/_00976_ ),
    .Y(\soc/cpu/_02903_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07492_  (.A1(\soc/cpu/cpuregs_rdata2[1] ),
    .A2(\soc/cpu/_01414_ ),
    .B1(\soc/cpu/is_slli_srli_srai ),
    .Y(\soc/cpu/_02904_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/_07494_  (.A1(\soc/cpu/is_slli_srli_srai ),
    .A2(\soc/cpu/_02752_ ),
    .B1(\soc/cpu/_02904_ ),
    .C1(\soc/cpu/cpu_state[4] ),
    .X(\soc/cpu/_02906_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07495_  (.A(\soc/cpu/_00938_ ),
    .B(\soc/cpu/_02903_ ),
    .C(\soc/cpu/_02906_ ),
    .Y(\soc/cpu/_00669_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07498_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/decoded_imm[0] ),
    .B1(\soc/cpu/_01429_ ),
    .Y(\soc/cpu/_02909_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07499_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/decoded_imm[0] ),
    .B1(\soc/cpu/_02909_ ),
    .Y(\soc/cpu/_02910_ ));
 sky130_fd_sc_hd__or3_4 \soc/cpu/_07500_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/cpu_state[5] ),
    .C(\soc/cpu/cpu_state[4] ),
    .X(\soc/cpu/_02911_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07505_  (.A(\soc/cpu/cpuregs_rdata1[0] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02916_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_07506_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_02916_ ),
    .Y(\soc/cpu/_02917_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_07507_  (.A1(\soc/cpu/reg_next_pc[0] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_02917_ ),
    .Y(\soc/cpu/_02918_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_07508_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/cpu_state[4] ),
    .C(\soc/cpu/_00936_ ),
    .X(\soc/cpu/_02919_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07509_  (.A1(\soc/cpu/pcpi_rs1 [4]),
    .A2(\soc/cpu/_01421_ ),
    .B1(\soc/cpu/_02919_ ),
    .Y(\soc/cpu/_02920_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_07510_  (.A1(\soc/cpu/_02911_ ),
    .A2(\soc/cpu/_02918_ ),
    .B1(\soc/cpu/_02920_ ),
    .B2(\soc/cpu/_02705_ ),
    .Y(\soc/cpu/_02921_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07511_  (.A1(\soc/cpu/_02910_ ),
    .A2(\soc/cpu/_02921_ ),
    .B1(net50),
    .Y(\soc/cpu/_02922_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07512_  (.A1(\soc/cpu/_01490_ ),
    .A2(net50),
    .B1(\soc/cpu/_02922_ ),
    .Y(\soc/cpu/_00670_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07514_  (.A(\soc/cpu/_02642_ ),
    .B(\soc/cpu/_02643_ ),
    .Y(\soc/cpu/_02924_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07515_  (.A(\soc/cpu/_02642_ ),
    .B(\soc/cpu/_02643_ ),
    .Y(\soc/cpu/_02925_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07516_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_02925_ ),
    .Y(\soc/cpu/_02926_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07517_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/_02705_ ),
    .Y(\soc/cpu/_02927_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07519_  (.A(\soc/cpu/pcpi_rs1 [0]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_02929_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07520_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_02927_ ),
    .C(\soc/cpu/_02929_ ),
    .Y(\soc/cpu/_02930_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07521_  (.A1(\soc/cpu/_02924_ ),
    .A2(\soc/cpu/_02926_ ),
    .B1(\soc/cpu/_02930_ ),
    .Y(\soc/cpu/_02931_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_07525_  (.A(\soc/cpu/cpuregs_rdata1[1] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02935_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07527_  (.A(\soc/cpu/reg_pc[1] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_02937_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07528_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_02935_ ),
    .B1(\soc/cpu/_02937_ ),
    .Y(\soc/cpu/_02938_ ));
 sky130_fd_sc_hd__a32oi_4 \soc/cpu/_07530_  (.A1(\soc/cpu/pcpi_rs1 [5]),
    .A2(\soc/cpu/_01421_ ),
    .A3(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_02938_ ),
    .B2(\soc/cpu/_02692_ ),
    .Y(\soc/cpu/_02940_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07532_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(net50),
    .Y(\soc/cpu/_02942_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07533_  (.A1(net50),
    .A2(\soc/cpu/_02931_ ),
    .A3(\soc/cpu/_02940_ ),
    .B1(\soc/cpu/_02942_ ),
    .Y(\soc/cpu/_00671_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07535_  (.A(\soc/cpu/_02641_ ),
    .B(\soc/cpu/_02645_ ),
    .X(\soc/cpu/_02944_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07536_  (.A(\soc/cpu/cpuregs_rdata1[2] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02945_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07537_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_02945_ ),
    .Y(\soc/cpu/_02946_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_07538_  (.A1(\soc/cpu/reg_pc[2] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_02946_ ),
    .Y(\soc/cpu/_02947_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07540_  (.A(\soc/cpu/pcpi_rs1 [1]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_02949_ ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_07541_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/_00936_ ),
    .X(\soc/cpu/_02950_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07542_  (.A1(\soc/cpu/pcpi_rs1 [3]),
    .A2(net156),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_02951_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07543_  (.A(\soc/cpu/_02949_ ),
    .B(\soc/cpu/_02951_ ),
    .Y(\soc/cpu/_02952_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07544_  (.A1(\soc/cpu/pcpi_rs1 [6]),
    .A2(\soc/cpu/_01421_ ),
    .A3(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_02952_ ),
    .Y(\soc/cpu/_02953_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07545_  (.A1(\soc/cpu/_02911_ ),
    .A2(\soc/cpu/_02947_ ),
    .B1(\soc/cpu/_02953_ ),
    .Y(\soc/cpu/_02954_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07546_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_02944_ ),
    .B1(\soc/cpu/_02954_ ),
    .Y(\soc/cpu/_02955_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07548_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(net50),
    .Y(\soc/cpu/_02957_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07549_  (.A1(net50),
    .A2(\soc/cpu/_02955_ ),
    .B1(\soc/cpu/_02957_ ),
    .Y(\soc/cpu/_00672_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07550_  (.A1(\soc/cpu/_02641_ ),
    .A2(\soc/cpu/_02645_ ),
    .B1(\soc/cpu/_02639_ ),
    .Y(\soc/cpu/_02958_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07551_  (.A(\soc/cpu/_02646_ ),
    .B(\soc/cpu/_02638_ ),
    .Y(\soc/cpu/_02959_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07552_  (.A(\soc/cpu/_02958_ ),
    .B(\soc/cpu/_02959_ ),
    .Y(\soc/cpu/_02960_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07553_  (.A(\soc/cpu/cpuregs_rdata1[3] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02961_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07554_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_02961_ ),
    .Y(\soc/cpu/_02962_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_07555_  (.A1(\soc/cpu/reg_pc[3] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_02962_ ),
    .Y(\soc/cpu/_02963_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07556_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/_02705_ ),
    .Y(\soc/cpu/_02964_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07557_  (.A(\soc/cpu/pcpi_rs1 [2]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_02965_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07558_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_02964_ ),
    .C(\soc/cpu/_02965_ ),
    .Y(\soc/cpu/_02966_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07559_  (.A1(\soc/cpu/pcpi_rs1 [7]),
    .A2(\soc/cpu/_01421_ ),
    .A3(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_02966_ ),
    .Y(\soc/cpu/_02967_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07560_  (.A1(\soc/cpu/_02911_ ),
    .A2(\soc/cpu/_02963_ ),
    .B1(\soc/cpu/_02967_ ),
    .Y(\soc/cpu/_02968_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07561_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_02960_ ),
    .B1(\soc/cpu/_02968_ ),
    .Y(\soc/cpu/_02969_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07562_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(net50),
    .Y(\soc/cpu/_02970_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07563_  (.A1(net50),
    .A2(\soc/cpu/_02969_ ),
    .B1(\soc/cpu/_02970_ ),
    .Y(\soc/cpu/_00673_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07564_  (.A1(\soc/cpu/_02638_ ),
    .A2(\soc/cpu/_02647_ ),
    .B1(\soc/cpu/_02637_ ),
    .Y(\soc/cpu/_02971_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07565_  (.A(\soc/cpu/_02637_ ),
    .B(\soc/cpu/_02638_ ),
    .C(\soc/cpu/_02647_ ),
    .Y(\soc/cpu/_02972_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07566_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_02972_ ),
    .Y(\soc/cpu/_02973_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07568_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(\soc/cpu/_02705_ ),
    .Y(\soc/cpu/_02975_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07569_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_02929_ ),
    .C(\soc/cpu/_02975_ ),
    .Y(\soc/cpu/_02976_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07571_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(net156),
    .Y(\soc/cpu/_02978_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07572_  (.A(\soc/cpu/pcpi_rs1 [3]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_02979_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_07573_  (.A(\soc/cpu/cpuregs_rdata1[4] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02980_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07574_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_02980_ ),
    .Y(\soc/cpu/_02981_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_07575_  (.A1(\soc/cpu/reg_pc[4] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_02981_ ),
    .Y(\soc/cpu/_02982_ ));
 sky130_fd_sc_hd__o32ai_4 \soc/cpu/_07576_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_02978_ ),
    .A3(\soc/cpu/_02979_ ),
    .B1(\soc/cpu/_02911_ ),
    .B2(\soc/cpu/_02982_ ),
    .Y(\soc/cpu/_02983_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07577_  (.A1(\soc/cpu/_02971_ ),
    .A2(\soc/cpu/_02973_ ),
    .B1(\soc/cpu/_02976_ ),
    .C1(\soc/cpu/_02983_ ),
    .Y(\soc/cpu/_02984_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07578_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(net50),
    .Y(\soc/cpu/_02985_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07579_  (.A1(net50),
    .A2(\soc/cpu/_02984_ ),
    .B1(\soc/cpu/_02985_ ),
    .Y(\soc/cpu/_00674_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07581_  (.A(\soc/cpu/cpuregs_rdata1[5] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_02987_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07582_  (.A(\soc/cpu/reg_pc[5] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_02988_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07583_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_02987_ ),
    .B1(\soc/cpu/_02988_ ),
    .Y(\soc/cpu/_02989_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07585_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(net156),
    .Y(\soc/cpu/_02991_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07586_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_02949_ ),
    .C(\soc/cpu/_02991_ ),
    .Y(\soc/cpu/_02992_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07587_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_02989_ ),
    .B1(\soc/cpu/_02992_ ),
    .Y(\soc/cpu/_02993_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07588_  (.A1(\soc/cpu/decoded_imm[4] ),
    .A2(\soc/cpu/pcpi_rs1 [4]),
    .B1(\soc/cpu/_02972_ ),
    .Y(\soc/cpu/_02994_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_07589_  (.A(\soc/cpu/_02649_ ),
    .SLEEP(\soc/cpu/_02636_ ),
    .X(\soc/cpu/_02995_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07590_  (.A(\soc/cpu/_02994_ ),
    .B(\soc/cpu/_02995_ ),
    .Y(\soc/cpu/_02996_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07591_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(\soc/cpu/_02705_ ),
    .Y(\soc/cpu/_02997_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07592_  (.A(\soc/cpu/pcpi_rs1 [4]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_02998_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07593_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_02997_ ),
    .C(\soc/cpu/_02998_ ),
    .Y(\soc/cpu/_02999_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07594_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_02996_ ),
    .B1(\soc/cpu/_02999_ ),
    .Y(\soc/cpu/_03000_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07595_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(net50),
    .Y(\soc/cpu/_03001_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07596_  (.A1(net50),
    .A2(\soc/cpu/_02993_ ),
    .A3(\soc/cpu/_03000_ ),
    .B1(\soc/cpu/_03001_ ),
    .Y(\soc/cpu/_00675_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07597_  (.A(\soc/cpu/_02636_ ),
    .B(\soc/cpu/_02650_ ),
    .Y(\soc/cpu/_03002_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07598_  (.A(\soc/cpu/_02635_ ),
    .B(\soc/cpu/_03002_ ),
    .Y(\soc/cpu/_03003_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07599_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(\soc/cpu/_02705_ ),
    .Y(\soc/cpu/_03004_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07600_  (.A(\soc/cpu/pcpi_rs1 [5]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03005_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07601_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_03004_ ),
    .C(\soc/cpu/_03005_ ),
    .Y(\soc/cpu/_03006_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07602_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(net156),
    .Y(\soc/cpu/_03007_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_07603_  (.A(\soc/cpu/cpuregs_rdata1[6] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03008_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07604_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03008_ ),
    .Y(\soc/cpu/_03009_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07605_  (.A1(\soc/cpu/reg_pc[6] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03009_ ),
    .Y(\soc/cpu/_03010_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07606_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_02965_ ),
    .A3(\soc/cpu/_03007_ ),
    .B1(\soc/cpu/_03010_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03011_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07607_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03003_ ),
    .B1(\soc/cpu/_03006_ ),
    .C1(\soc/cpu/_03011_ ),
    .Y(\soc/cpu/_03012_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07608_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(net50),
    .Y(\soc/cpu/_03013_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07609_  (.A1(net50),
    .A2(\soc/cpu/_03012_ ),
    .B1(\soc/cpu/_03013_ ),
    .Y(\soc/cpu/_00676_ ));
 sky130_fd_sc_hd__o31a_1 \soc/cpu/_07610_  (.A1(\soc/cpu/_02635_ ),
    .A2(\soc/cpu/_02636_ ),
    .A3(\soc/cpu/_02650_ ),
    .B1(\soc/cpu/_02651_ ),
    .X(\soc/cpu/_03014_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_07611_  (.A(\soc/cpu/_02652_ ),
    .SLEEP(\soc/cpu/_02634_ ),
    .X(\soc/cpu/_03015_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07612_  (.A(\soc/cpu/_03014_ ),
    .B(\soc/cpu/_03015_ ),
    .Y(\soc/cpu/_03016_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07613_  (.A(\soc/cpu/pcpi_rs1 [6]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03017_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07614_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_02975_ ),
    .C(\soc/cpu/_03017_ ),
    .Y(\soc/cpu/_03018_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07615_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(net156),
    .Y(\soc/cpu/_03019_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_07617_  (.A(\soc/cpu/cpuregs_rdata1[7] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03021_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07618_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03021_ ),
    .Y(\soc/cpu/_03022_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07619_  (.A1(\soc/cpu/reg_pc[7] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03022_ ),
    .Y(\soc/cpu/_03023_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07620_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_02979_ ),
    .A3(\soc/cpu/_03019_ ),
    .B1(\soc/cpu/_03023_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03024_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07621_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03016_ ),
    .B1(\soc/cpu/_03018_ ),
    .C1(\soc/cpu/_03024_ ),
    .Y(\soc/cpu/_03025_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07622_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(net49),
    .Y(\soc/cpu/_03026_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07623_  (.A1(net49),
    .A2(\soc/cpu/_03025_ ),
    .B1(\soc/cpu/_03026_ ),
    .Y(\soc/cpu/_00677_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07624_  (.A1(\soc/cpu/_02634_ ),
    .A2(\soc/cpu/_02653_ ),
    .B1(\soc/cpu/_02633_ ),
    .Y(\soc/cpu/_03027_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07625_  (.A(\soc/cpu/_02633_ ),
    .B(\soc/cpu/_02634_ ),
    .C(\soc/cpu/_02653_ ),
    .Y(\soc/cpu/_03028_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07626_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_03028_ ),
    .Y(\soc/cpu/_03029_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07627_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(net156),
    .Y(\soc/cpu/_03030_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07628_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_02998_ ),
    .C(\soc/cpu/_03030_ ),
    .Y(\soc/cpu/_03031_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07629_  (.A(\soc/cpu/pcpi_rs1 [7]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03032_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07630_  (.A(\soc/cpu/cpuregs_rdata1[8] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03033_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07631_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03033_ ),
    .Y(\soc/cpu/_03034_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07632_  (.A1(\soc/cpu/reg_pc[8] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03034_ ),
    .Y(\soc/cpu/_03035_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07633_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_02991_ ),
    .A3(\soc/cpu/_03032_ ),
    .B1(\soc/cpu/_03035_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03036_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07634_  (.A1(\soc/cpu/_03027_ ),
    .A2(\soc/cpu/_03029_ ),
    .B1(\soc/cpu/_03031_ ),
    .C1(\soc/cpu/_03036_ ),
    .Y(\soc/cpu/_03037_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07635_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(net49),
    .Y(\soc/cpu/_03038_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07636_  (.A1(net49),
    .A2(\soc/cpu/_03037_ ),
    .B1(\soc/cpu/_03038_ ),
    .Y(\soc/cpu/_00678_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07637_  (.A1(\soc/cpu/decoded_imm[8] ),
    .A2(\soc/cpu/pcpi_rs1 [8]),
    .B1(\soc/cpu/_03028_ ),
    .Y(\soc/cpu/_03039_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07638_  (.A(\soc/cpu/_02655_ ),
    .B(\soc/cpu/_02632_ ),
    .Y(\soc/cpu/_03040_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07639_  (.A(\soc/cpu/_03039_ ),
    .B(\soc/cpu/_03040_ ),
    .X(\soc/cpu/_03041_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07640_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(net156),
    .Y(\soc/cpu/_03042_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07641_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_03005_ ),
    .C(\soc/cpu/_03042_ ),
    .Y(\soc/cpu/_03043_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07642_  (.A(\soc/cpu/pcpi_rs1 [8]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03044_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07643_  (.A(\soc/cpu/cpuregs_rdata1[9] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03045_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07644_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03045_ ),
    .Y(\soc/cpu/_03046_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07645_  (.A1(\soc/cpu/reg_pc[9] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03046_ ),
    .Y(\soc/cpu/_03047_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07646_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03007_ ),
    .A3(\soc/cpu/_03044_ ),
    .B1(\soc/cpu/_03047_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03048_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07647_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03041_ ),
    .B1(\soc/cpu/_03043_ ),
    .C1(\soc/cpu/_03048_ ),
    .Y(\soc/cpu/_03049_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07648_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(net49),
    .Y(\soc/cpu/_03050_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07649_  (.A1(net49),
    .A2(\soc/cpu/_03049_ ),
    .B1(\soc/cpu/_03050_ ),
    .Y(\soc/cpu/_00679_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07650_  (.A(\soc/cpu/_02632_ ),
    .B(\soc/cpu/_02656_ ),
    .X(\soc/cpu/_03051_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07651_  (.A1(\soc/cpu/_02631_ ),
    .A2(\soc/cpu/_03051_ ),
    .B1(\soc/cpu/_01429_ ),
    .Y(\soc/cpu/_03052_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07652_  (.A1(\soc/cpu/_02631_ ),
    .A2(\soc/cpu/_03051_ ),
    .B1(\soc/cpu/_03052_ ),
    .Y(\soc/cpu/_03053_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07653_  (.A(\soc/cpu/pcpi_rs1 [9]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03054_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07654_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_03019_ ),
    .C(\soc/cpu/_03054_ ),
    .Y(\soc/cpu/_03055_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07655_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(net156),
    .Y(\soc/cpu/_03056_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07656_  (.A(\soc/cpu/cpuregs_rdata1[10] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03057_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07657_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03057_ ),
    .Y(\soc/cpu/_03058_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07658_  (.A1(\soc/cpu/reg_pc[10] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03058_ ),
    .Y(\soc/cpu/_03059_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07659_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03017_ ),
    .A3(\soc/cpu/_03056_ ),
    .B1(\soc/cpu/_03059_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03060_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07660_  (.A1(\soc/cpu/_03053_ ),
    .A2(\soc/cpu/_03055_ ),
    .A3(\soc/cpu/_03060_ ),
    .B1(net49),
    .Y(\soc/cpu/_03061_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07661_  (.A1(\soc/cpu/_01535_ ),
    .A2(net50),
    .B1(\soc/cpu/_03061_ ),
    .Y(\soc/cpu/_00680_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07662_  (.A1(\soc/cpu/_02631_ ),
    .A2(\soc/cpu/_03051_ ),
    .B1(\soc/cpu/_02629_ ),
    .Y(\soc/cpu/_03062_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07663_  (.A(\soc/cpu/_02657_ ),
    .B(\soc/cpu/_02628_ ),
    .Y(\soc/cpu/_03063_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07664_  (.A(\soc/cpu/_03062_ ),
    .B(\soc/cpu/_03063_ ),
    .Y(\soc/cpu/_03064_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07665_  (.A(\soc/cpu/pcpi_rs1 [10]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03065_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07666_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_03030_ ),
    .C(\soc/cpu/_03065_ ),
    .Y(\soc/cpu/_03066_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07667_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(net156),
    .Y(\soc/cpu/_03067_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07668_  (.A(\soc/cpu/cpuregs_rdata1[11] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03068_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07669_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03068_ ),
    .Y(\soc/cpu/_03069_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07670_  (.A1(\soc/cpu/reg_pc[11] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03069_ ),
    .Y(\soc/cpu/_03070_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07671_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03032_ ),
    .A3(\soc/cpu/_03067_ ),
    .B1(\soc/cpu/_03070_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03071_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07672_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03064_ ),
    .B1(\soc/cpu/_03066_ ),
    .C1(\soc/cpu/_03071_ ),
    .Y(\soc/cpu/_03072_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07673_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(net49),
    .Y(\soc/cpu/_03073_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07674_  (.A1(net49),
    .A2(\soc/cpu/_03072_ ),
    .B1(\soc/cpu/_03073_ ),
    .Y(\soc/cpu/_00681_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07675_  (.A(\soc/cpu/_02627_ ),
    .B(\soc/cpu/_02628_ ),
    .C(\soc/cpu/_02658_ ),
    .Y(\soc/cpu/_03074_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_07676_  (.A1(\soc/cpu/_02628_ ),
    .A2(\soc/cpu/_02658_ ),
    .B1(\soc/cpu/_02627_ ),
    .X(\soc/cpu/_03075_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07677_  (.A(\soc/cpu/cpuregs_rdata1[12] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03076_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07678_  (.A(\soc/cpu/reg_pc[12] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03077_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07679_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03076_ ),
    .B1(\soc/cpu/_03077_ ),
    .Y(\soc/cpu/_03078_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07680_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(net156),
    .Y(\soc/cpu/_03079_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07681_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_03044_ ),
    .C(\soc/cpu/_03079_ ),
    .Y(\soc/cpu/_03080_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07682_  (.A(\soc/cpu/pcpi_rs1 [11]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03081_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07683_  (.A(\soc/cpu/_00937_ ),
    .B(\soc/cpu/_03042_ ),
    .C(\soc/cpu/_03081_ ),
    .Y(\soc/cpu/_03082_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07684_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03078_ ),
    .B1(\soc/cpu/_03080_ ),
    .C1(\soc/cpu/_03082_ ),
    .Y(\soc/cpu/_03083_ ));
 sky130_fd_sc_hd__o311ai_1 \soc/cpu/_07685_  (.A1(\soc/cpu/_00838_ ),
    .A2(\soc/cpu/_03074_ ),
    .A3(\soc/cpu/_03075_ ),
    .B1(\soc/cpu/_03083_ ),
    .C1(net49),
    .Y(\soc/cpu/_03084_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_07686_  (.A1(\soc/cpu/pcpi_rs1 [12]),
    .A2(net49),
    .B1(\soc/cpu/_03084_ ),
    .X(\soc/cpu/_00682_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07687_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(net49),
    .Y(\soc/cpu/_03085_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07688_  (.A1(\soc/cpu/decoded_imm[12] ),
    .A2(\soc/cpu/pcpi_rs1 [12]),
    .B1(\soc/cpu/_03074_ ),
    .Y(\soc/cpu/_03086_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07689_  (.A(\soc/cpu/_02660_ ),
    .B(\soc/cpu/_02626_ ),
    .Y(\soc/cpu/_03087_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07690_  (.A(\soc/cpu/_03086_ ),
    .B(\soc/cpu/_03087_ ),
    .X(\soc/cpu/_03088_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07691_  (.A(\soc/cpu/pcpi_rs1 [12]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03089_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07692_  (.A(\soc/cpu/cpuregs_rdata1[13] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03090_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07693_  (.A(\soc/cpu/reg_pc[13] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03091_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07694_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03090_ ),
    .B1(\soc/cpu/_03091_ ),
    .Y(\soc/cpu/_03092_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07695_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(net156),
    .Y(\soc/cpu/_03093_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07696_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_03054_ ),
    .C(\soc/cpu/_03093_ ),
    .Y(\soc/cpu/_03094_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07697_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03092_ ),
    .B1(\soc/cpu/_03094_ ),
    .Y(\soc/cpu/_03095_ ));
 sky130_fd_sc_hd__o311ai_2 \soc/cpu/_07698_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03056_ ),
    .A3(\soc/cpu/_03089_ ),
    .B1(\soc/cpu/_03095_ ),
    .C1(net49),
    .Y(\soc/cpu/_03096_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07699_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03088_ ),
    .B1(\soc/cpu/_03096_ ),
    .Y(\soc/cpu/_03097_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07700_  (.A(\soc/cpu/_03085_ ),
    .B(\soc/cpu/_03097_ ),
    .Y(\soc/cpu/_00683_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_07701_  (.A(\soc/cpu/_02626_ ),
    .B(\soc/cpu/_02661_ ),
    .X(\soc/cpu/_03098_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_07702_  (.A(\soc/cpu/_02625_ ),
    .B(\soc/cpu/_02626_ ),
    .C(\soc/cpu/_02661_ ),
    .X(\soc/cpu/_03099_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07703_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_03099_ ),
    .Y(\soc/cpu/_03100_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07704_  (.A1(\soc/cpu/_02625_ ),
    .A2(\soc/cpu/_03098_ ),
    .B1(\soc/cpu/_03100_ ),
    .Y(\soc/cpu/_03101_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07705_  (.A(\soc/cpu/cpuregs_rdata1[14] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03102_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07706_  (.A(\soc/cpu/reg_pc[14] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03103_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07707_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03102_ ),
    .B1(\soc/cpu/_03103_ ),
    .Y(\soc/cpu/_03104_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07708_  (.A(\soc/cpu/pcpi_rs1 [13]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03105_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07709_  (.A1(\soc/cpu/pcpi_rs1 [18]),
    .A2(net156),
    .B1(\soc/cpu/_01421_ ),
    .Y(\soc/cpu/_03106_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07710_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03067_ ),
    .A3(\soc/cpu/_03105_ ),
    .B1(\soc/cpu/_03106_ ),
    .B2(\soc/cpu/_03065_ ),
    .Y(\soc/cpu/_03107_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07711_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03104_ ),
    .B1(\soc/cpu/_03107_ ),
    .Y(\soc/cpu/_03108_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07712_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(net49),
    .Y(\soc/cpu/_03109_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07713_  (.A1(net49),
    .A2(\soc/cpu/_03101_ ),
    .A3(\soc/cpu/_03108_ ),
    .B1(\soc/cpu/_03109_ ),
    .Y(\soc/cpu/_00684_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07714_  (.A(\soc/cpu/_02623_ ),
    .B(\soc/cpu/_03099_ ),
    .Y(\soc/cpu/_03110_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07715_  (.A(\soc/cpu/_02622_ ),
    .B(\soc/cpu/_02662_ ),
    .Y(\soc/cpu/_03111_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07716_  (.A(\soc/cpu/_03110_ ),
    .B(\soc/cpu/_03111_ ),
    .Y(\soc/cpu/_03112_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07717_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(net156),
    .Y(\soc/cpu/_03113_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07718_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_03081_ ),
    .C(\soc/cpu/_03113_ ),
    .Y(\soc/cpu/_03114_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07719_  (.A(\soc/cpu/pcpi_rs1 [14]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03115_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07720_  (.A(\soc/cpu/cpuregs_rdata1[15] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03116_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07721_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03116_ ),
    .Y(\soc/cpu/_03117_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07722_  (.A1(\soc/cpu/reg_pc[15] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03117_ ),
    .Y(\soc/cpu/_03118_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07723_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03079_ ),
    .A3(\soc/cpu/_03115_ ),
    .B1(\soc/cpu/_03118_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03119_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07724_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03112_ ),
    .B1(\soc/cpu/_03114_ ),
    .C1(\soc/cpu/_03119_ ),
    .Y(\soc/cpu/_03120_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07725_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(net48),
    .Y(\soc/cpu/_03121_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07726_  (.A1(net49),
    .A2(\soc/cpu/_03120_ ),
    .B1(\soc/cpu/_03121_ ),
    .Y(\soc/cpu/_00685_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07727_  (.A(\soc/cpu/_02622_ ),
    .B(\soc/cpu/_02663_ ),
    .Y(\soc/cpu/_03122_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07728_  (.A(\soc/cpu/_02621_ ),
    .B(\soc/cpu/_03122_ ),
    .X(\soc/cpu/_03123_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07729_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_03123_ ),
    .Y(\soc/cpu/_03124_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07730_  (.A(\soc/cpu/pcpi_rs1 [15]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03125_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07731_  (.A(\soc/cpu/cpuregs_rdata1[16] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03126_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07732_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03126_ ),
    .Y(\soc/cpu/_03127_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07733_  (.A1(\soc/cpu/reg_pc[16] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03127_ ),
    .Y(\soc/cpu/_03128_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07734_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03093_ ),
    .A3(\soc/cpu/_03125_ ),
    .B1(\soc/cpu/_03128_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03129_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07735_  (.A1(\soc/cpu/pcpi_rs1 [20]),
    .A2(net156),
    .B1(\soc/cpu/_01421_ ),
    .Y(\soc/cpu/_03130_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07736_  (.A1(\soc/cpu/_03089_ ),
    .A2(\soc/cpu/_03130_ ),
    .B1(net48),
    .Y(\soc/cpu/_03131_ ));
 sky130_fd_sc_hd__o32a_1 \soc/cpu/_07737_  (.A1(\soc/cpu/_03124_ ),
    .A2(\soc/cpu/_03129_ ),
    .A3(\soc/cpu/_03131_ ),
    .B1(net48),
    .B2(\soc/cpu/pcpi_rs1 [16]),
    .X(\soc/cpu/_00686_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07738_  (.A1(\soc/cpu/_02621_ ),
    .A2(\soc/cpu/_02622_ ),
    .A3(\soc/cpu/_02663_ ),
    .B1(\soc/cpu/_02664_ ),
    .Y(\soc/cpu/_03132_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07739_  (.A(\soc/cpu/_02665_ ),
    .B(\soc/cpu/_02620_ ),
    .Y(\soc/cpu/_03133_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07740_  (.A(\soc/cpu/_03132_ ),
    .B(\soc/cpu/_03133_ ),
    .Y(\soc/cpu/_03134_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07742_  (.A(\soc/cpu/cpuregs_rdata1[17] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03136_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07743_  (.A(\soc/cpu/reg_pc[17] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03137_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07744_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03136_ ),
    .B1(\soc/cpu/_03137_ ),
    .Y(\soc/cpu/_03138_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07745_  (.A(\soc/cpu/pcpi_rs1 [21]),
    .B(net155),
    .Y(\soc/cpu/_03139_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07746_  (.A1(\soc/cpu/pcpi_rs1 [18]),
    .A2(net155),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03140_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07747_  (.A(\soc/cpu/pcpi_rs1 [16]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03141_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07748_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03105_ ),
    .A3(\soc/cpu/_03139_ ),
    .B1(\soc/cpu/_03140_ ),
    .B2(\soc/cpu/_03141_ ),
    .Y(\soc/cpu/_03142_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07749_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03134_ ),
    .B1(\soc/cpu/_03138_ ),
    .B2(\soc/cpu/_02692_ ),
    .C1(\soc/cpu/_03142_ ),
    .Y(\soc/cpu/_03143_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07750_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(net48),
    .Y(\soc/cpu/_03144_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07751_  (.A1(net48),
    .A2(\soc/cpu/_03143_ ),
    .B1(\soc/cpu/_03144_ ),
    .Y(\soc/cpu/_00687_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07752_  (.A1(\soc/cpu/_02620_ ),
    .A2(\soc/cpu/_02666_ ),
    .B1(\soc/cpu/_02619_ ),
    .Y(\soc/cpu/_03145_ ));
 sky130_fd_sc_hd__a311oi_1 \soc/cpu/_07753_  (.A1(\soc/cpu/_02619_ ),
    .A2(\soc/cpu/_02620_ ),
    .A3(\soc/cpu/_02666_ ),
    .B1(\soc/cpu/_03145_ ),
    .C1(\soc/cpu/_00838_ ),
    .Y(\soc/cpu/_03146_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07754_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(net155),
    .Y(\soc/cpu/_03147_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07755_  (.A(\soc/cpu/cpuregs_rdata1[18] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03148_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07756_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03148_ ),
    .Y(\soc/cpu/_03149_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07757_  (.A1(\soc/cpu/reg_pc[18] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03149_ ),
    .Y(\soc/cpu/_03150_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07758_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03115_ ),
    .A3(\soc/cpu/_03147_ ),
    .B1(\soc/cpu/_03150_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03151_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07759_  (.A(\soc/cpu/pcpi_rs1 [17]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03152_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07760_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03113_ ),
    .A3(\soc/cpu/_03152_ ),
    .B1(net48),
    .Y(\soc/cpu/_03153_ ));
 sky130_fd_sc_hd__o32a_1 \soc/cpu/_07761_  (.A1(\soc/cpu/_03146_ ),
    .A2(\soc/cpu/_03151_ ),
    .A3(\soc/cpu/_03153_ ),
    .B1(net48),
    .B2(\soc/cpu/pcpi_rs1 [18]),
    .X(\soc/cpu/_00688_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_07762_  (.A(\soc/cpu/_02616_ ),
    .SLEEP(\soc/cpu/_02668_ ),
    .X(\soc/cpu/_03154_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07763_  (.A(\soc/cpu/_02667_ ),
    .B(\soc/cpu/_03154_ ),
    .Y(\soc/cpu/_03155_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07764_  (.A(\soc/cpu/_01429_ ),
    .B(\soc/cpu/_03155_ ),
    .Y(\soc/cpu/_03156_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07765_  (.A(\soc/cpu/cpuregs_rdata1[19] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03157_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07766_  (.A(\soc/cpu/reg_pc[19] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03158_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_07767_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03157_ ),
    .B1(\soc/cpu/_03158_ ),
    .Y(\soc/cpu/_03159_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07768_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(net155),
    .Y(\soc/cpu/_03160_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07769_  (.A(\soc/cpu/pcpi_rs1 [18]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03161_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07770_  (.A1(\soc/cpu/pcpi_rs1 [20]),
    .A2(net155),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03162_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07771_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03125_ ),
    .A3(\soc/cpu/_03160_ ),
    .B1(\soc/cpu/_03161_ ),
    .B2(\soc/cpu/_03162_ ),
    .Y(\soc/cpu/_03163_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07772_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03159_ ),
    .B1(\soc/cpu/_03163_ ),
    .Y(\soc/cpu/_03164_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07773_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(net48),
    .Y(\soc/cpu/_03165_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07774_  (.A1(net48),
    .A2(\soc/cpu/_03156_ ),
    .A3(\soc/cpu/_03164_ ),
    .B1(\soc/cpu/_03165_ ),
    .Y(\soc/cpu/_00689_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07775_  (.A(\soc/cpu/decoded_imm[20] ),
    .B(\soc/cpu/pcpi_rs1 [20]),
    .X(\soc/cpu/_03166_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07776_  (.A(\soc/cpu/_03166_ ),
    .B(\soc/cpu/_02669_ ),
    .Y(\soc/cpu/_03167_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07777_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_03167_ ),
    .Y(\soc/cpu/_03168_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07778_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(net155),
    .Y(\soc/cpu/_03169_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07779_  (.A(\soc/cpu/cpuregs_rdata1[20] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03170_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07780_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03170_ ),
    .Y(\soc/cpu/_03171_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_07781_  (.A1(\soc/cpu/reg_pc[20] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03171_ ),
    .Y(\soc/cpu/_03172_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07782_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03141_ ),
    .A3(\soc/cpu/_03169_ ),
    .B1(\soc/cpu/_03172_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03173_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07783_  (.A(\soc/cpu/pcpi_rs1 [19]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03174_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07784_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03139_ ),
    .A3(\soc/cpu/_03174_ ),
    .B1(net48),
    .Y(\soc/cpu/_03175_ ));
 sky130_fd_sc_hd__o32a_1 \soc/cpu/_07785_  (.A1(\soc/cpu/_03168_ ),
    .A2(\soc/cpu/_03173_ ),
    .A3(\soc/cpu/_03175_ ),
    .B1(net48),
    .B2(\soc/cpu/pcpi_rs1 [20]),
    .X(\soc/cpu/_00690_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07786_  (.A(\soc/cpu/decoded_imm[21] ),
    .B(\soc/cpu/pcpi_rs1 [21]),
    .X(\soc/cpu/_03176_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07787_  (.A(\soc/cpu/_02670_ ),
    .B(\soc/cpu/_03176_ ),
    .Y(\soc/cpu/_03177_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07788_  (.A(\soc/cpu/_00838_ ),
    .B(\soc/cpu/_03177_ ),
    .Y(\soc/cpu/_03178_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07789_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .B(net155),
    .Y(\soc/cpu/_03179_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07790_  (.A(\soc/cpu/cpuregs_rdata1[21] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03180_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07791_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03180_ ),
    .Y(\soc/cpu/_03181_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_07792_  (.A1(\soc/cpu/reg_pc[21] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03181_ ),
    .Y(\soc/cpu/_03182_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07793_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03152_ ),
    .A3(\soc/cpu/_03179_ ),
    .B1(\soc/cpu/_03182_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03183_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07794_  (.A(\soc/cpu/pcpi_rs1 [20]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03184_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07795_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03147_ ),
    .A3(\soc/cpu/_03184_ ),
    .B1(net48),
    .Y(\soc/cpu/_03185_ ));
 sky130_fd_sc_hd__o32a_1 \soc/cpu/_07796_  (.A1(\soc/cpu/_03178_ ),
    .A2(\soc/cpu/_03183_ ),
    .A3(\soc/cpu/_03185_ ),
    .B1(net48),
    .B2(\soc/cpu/pcpi_rs1 [21]),
    .X(\soc/cpu/_00691_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_07797_  (.A_N(\soc/cpu/_02672_ ),
    .B(\soc/cpu/_02615_ ),
    .Y(\soc/cpu/_03186_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07798_  (.A(\soc/cpu/_03186_ ),
    .B(\soc/cpu/_02671_ ),
    .Y(\soc/cpu/_03187_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07799_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(net155),
    .Y(\soc/cpu/_03188_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07800_  (.A(\soc/cpu/_01409_ ),
    .B(\soc/cpu/_03161_ ),
    .C(\soc/cpu/_03188_ ),
    .Y(\soc/cpu/_03189_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07801_  (.A(\soc/cpu/pcpi_rs1 [21]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03190_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07802_  (.A(\soc/cpu/cpuregs_rdata1[22] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03191_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07803_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03191_ ),
    .Y(\soc/cpu/_03192_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07804_  (.A1(\soc/cpu/reg_pc[22] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03192_ ),
    .Y(\soc/cpu/_03193_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/cpu/_07805_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03160_ ),
    .A3(\soc/cpu/_03190_ ),
    .B1(\soc/cpu/_03193_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03194_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07806_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03187_ ),
    .B1(\soc/cpu/_03189_ ),
    .C1(\soc/cpu/_03194_ ),
    .Y(\soc/cpu/_03195_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07807_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(net48),
    .Y(\soc/cpu/_03196_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07808_  (.A1(net48),
    .A2(\soc/cpu/_03195_ ),
    .B1(\soc/cpu/_03196_ ),
    .Y(\soc/cpu/_00692_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_07809_  (.A(\soc/cpu/_02614_ ),
    .SLEEP(\soc/cpu/_02674_ ),
    .X(\soc/cpu/_03197_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07810_  (.A(\soc/cpu/_02673_ ),
    .B(\soc/cpu/_03197_ ),
    .Y(\soc/cpu/_03198_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07811_  (.A(\soc/cpu/_01429_ ),
    .B(\soc/cpu/_03198_ ),
    .Y(\soc/cpu/_03199_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07812_  (.A(\soc/cpu/cpuregs_rdata1[23] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03200_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07813_  (.A(\soc/cpu/reg_pc[23] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03201_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07814_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03200_ ),
    .B1(\soc/cpu/_03201_ ),
    .Y(\soc/cpu/_03202_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07815_  (.A(\soc/cpu/pcpi_rs1 [22]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03203_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07816_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(net155),
    .B1(\soc/cpu/_01421_ ),
    .Y(\soc/cpu/_03204_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07817_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03169_ ),
    .A3(\soc/cpu/_03203_ ),
    .B1(\soc/cpu/_03204_ ),
    .B2(\soc/cpu/_03174_ ),
    .Y(\soc/cpu/_03205_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07818_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03202_ ),
    .B1(\soc/cpu/_03205_ ),
    .Y(\soc/cpu/_03206_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07819_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(net47),
    .Y(\soc/cpu/_03207_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07820_  (.A1(net47),
    .A2(\soc/cpu/_03199_ ),
    .A3(\soc/cpu/_03206_ ),
    .B1(\soc/cpu/_03207_ ),
    .Y(\soc/cpu/_00693_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07821_  (.A1(\soc/cpu/_02614_ ),
    .A2(\soc/cpu/_02673_ ),
    .B1(\soc/cpu/_02674_ ),
    .Y(\soc/cpu/_03208_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07822_  (.A(\soc/cpu/_02675_ ),
    .B(\soc/cpu/_03208_ ),
    .Y(\soc/cpu/_03209_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07823_  (.A(\soc/cpu/_01429_ ),
    .B(\soc/cpu/_03209_ ),
    .Y(\soc/cpu/_03210_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07824_  (.A(\soc/cpu/cpuregs_rdata1[24] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03211_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07825_  (.A(\soc/cpu/reg_pc[24] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03212_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07826_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03211_ ),
    .B1(\soc/cpu/_03212_ ),
    .Y(\soc/cpu/_03213_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07827_  (.A(\soc/cpu/pcpi_rs1 [23]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03214_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07828_  (.A1(\soc/cpu/pcpi_rs1 [28]),
    .A2(net155),
    .B1(\soc/cpu/_01421_ ),
    .Y(\soc/cpu/_03215_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07829_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03179_ ),
    .A3(\soc/cpu/_03214_ ),
    .B1(\soc/cpu/_03215_ ),
    .B2(\soc/cpu/_03184_ ),
    .Y(\soc/cpu/_03216_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07830_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03213_ ),
    .B1(\soc/cpu/_03216_ ),
    .Y(\soc/cpu/_03217_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07831_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(net47),
    .Y(\soc/cpu/_03218_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07832_  (.A1(net47),
    .A2(\soc/cpu/_03210_ ),
    .A3(\soc/cpu/_03217_ ),
    .B1(\soc/cpu/_03218_ ),
    .Y(\soc/cpu/_00694_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07833_  (.A(\soc/cpu/decoded_imm[25] ),
    .B(\soc/cpu/pcpi_rs1 [25]),
    .Y(\soc/cpu/_03219_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07834_  (.A1(\soc/cpu/_02677_ ),
    .A2(\soc/cpu/_03219_ ),
    .B1(\soc/cpu/_01429_ ),
    .Y(\soc/cpu/_03220_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07835_  (.A1(\soc/cpu/_02677_ ),
    .A2(\soc/cpu/_03219_ ),
    .B1(\soc/cpu/_03220_ ),
    .Y(\soc/cpu/_03221_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07836_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(net155),
    .Y(\soc/cpu/_03222_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07837_  (.A(\soc/cpu/cpuregs_rdata1[25] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03223_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07838_  (.A(\soc/cpu/is_lui_auipc_jal ),
    .B(\soc/cpu/_03223_ ),
    .Y(\soc/cpu/_03224_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07839_  (.A1(\soc/cpu/reg_pc[25] ),
    .A2(\soc/cpu/_02699_ ),
    .B1(\soc/cpu/_03224_ ),
    .Y(\soc/cpu/_03225_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07840_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03190_ ),
    .A3(\soc/cpu/_03222_ ),
    .B1(\soc/cpu/_03225_ ),
    .B2(\soc/cpu/_02911_ ),
    .Y(\soc/cpu/_03226_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07841_  (.A(\soc/cpu/pcpi_rs1 [24]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03227_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07842_  (.A1(\soc/cpu/_00937_ ),
    .A2(\soc/cpu/_03188_ ),
    .A3(\soc/cpu/_03227_ ),
    .B1(net48),
    .Y(\soc/cpu/_03228_ ));
 sky130_fd_sc_hd__o32a_1 \soc/cpu/_07843_  (.A1(\soc/cpu/_03221_ ),
    .A2(\soc/cpu/_03226_ ),
    .A3(\soc/cpu/_03228_ ),
    .B1(net47),
    .B2(\soc/cpu/pcpi_rs1 [25]),
    .X(\soc/cpu/_00695_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07844_  (.A1(\soc/cpu/_02613_ ),
    .A2(\soc/cpu/_02677_ ),
    .B1(\soc/cpu/_02678_ ),
    .Y(\soc/cpu/_03229_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07845_  (.A(\soc/cpu/_02679_ ),
    .B(\soc/cpu/_03229_ ),
    .Y(\soc/cpu/_03230_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07846_  (.A(\soc/cpu/_01429_ ),
    .B(\soc/cpu/_03230_ ),
    .Y(\soc/cpu/_03231_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07847_  (.A(\soc/cpu/cpuregs_rdata1[26] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03232_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07848_  (.A(\soc/cpu/reg_pc[26] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03233_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07849_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03232_ ),
    .B1(\soc/cpu/_03233_ ),
    .Y(\soc/cpu/_03234_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07850_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(net155),
    .Y(\soc/cpu/_03235_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07851_  (.A(\soc/cpu/pcpi_rs1 [25]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03236_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07852_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(net155),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03237_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07853_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03203_ ),
    .A3(\soc/cpu/_03235_ ),
    .B1(\soc/cpu/_03236_ ),
    .B2(\soc/cpu/_03237_ ),
    .Y(\soc/cpu/_03238_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07854_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03234_ ),
    .B1(\soc/cpu/_03238_ ),
    .Y(\soc/cpu/_03239_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07855_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(net47),
    .Y(\soc/cpu/_03240_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07856_  (.A1(net47),
    .A2(\soc/cpu/_03231_ ),
    .A3(\soc/cpu/_03239_ ),
    .B1(\soc/cpu/_03240_ ),
    .Y(\soc/cpu/_00696_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_07857_  (.A(\soc/cpu/_02612_ ),
    .SLEEP(\soc/cpu/_02682_ ),
    .X(\soc/cpu/_03241_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_07858_  (.A(\soc/cpu/_02681_ ),
    .B(\soc/cpu/_03241_ ),
    .Y(\soc/cpu/_03242_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07859_  (.A(\soc/cpu/cpuregs_rdata1[27] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03243_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07860_  (.A(\soc/cpu/reg_pc[27] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03244_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07861_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03243_ ),
    .B1(\soc/cpu/_03244_ ),
    .Y(\soc/cpu/_03245_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07862_  (.A(\soc/cpu/pcpi_rs1 [31]),
    .B(net155),
    .Y(\soc/cpu/_03246_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07863_  (.A(\soc/cpu/pcpi_rs1 [26]),
    .B(\soc/cpu/_02603_ ),
    .Y(\soc/cpu/_03247_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07864_  (.A1(\soc/cpu/pcpi_rs1 [28]),
    .A2(net155),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03248_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/_07865_  (.A1(\soc/cpu/_01409_ ),
    .A2(\soc/cpu/_03214_ ),
    .A3(\soc/cpu/_03246_ ),
    .B1(\soc/cpu/_03247_ ),
    .B2(\soc/cpu/_03248_ ),
    .Y(\soc/cpu/_03249_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_07866_  (.A1(\soc/cpu/_01429_ ),
    .A2(\soc/cpu/_03242_ ),
    .B1(\soc/cpu/_03245_ ),
    .B2(\soc/cpu/_02692_ ),
    .C1(\soc/cpu/_03249_ ),
    .Y(\soc/cpu/_03250_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07867_  (.A(\soc/cpu/pcpi_rs1 [27]),
    .B(net47),
    .Y(\soc/cpu/_03251_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07868_  (.A1(net47),
    .A2(\soc/cpu/_03250_ ),
    .B1(\soc/cpu/_03251_ ),
    .Y(\soc/cpu/_00697_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_07869_  (.A(\soc/cpu/decoded_imm[28] ),
    .B(\soc/cpu/pcpi_rs1 [28]),
    .X(\soc/cpu/_03252_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07870_  (.A1(\soc/cpu/_03252_ ),
    .A2(\soc/cpu/_02683_ ),
    .B1(\soc/cpu/_00838_ ),
    .Y(\soc/cpu/_03253_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07871_  (.A1(\soc/cpu/_03252_ ),
    .A2(\soc/cpu/_02683_ ),
    .B1(\soc/cpu/_03253_ ),
    .Y(\soc/cpu/_03254_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07872_  (.A(\soc/cpu/cpuregs_rdata1[28] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03255_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07873_  (.A(\soc/cpu/reg_pc[28] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03256_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_07874_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03255_ ),
    .B1(\soc/cpu/_03256_ ),
    .Y(\soc/cpu/_03257_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07875_  (.A1(\soc/cpu/_02601_ ),
    .A2(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_03246_ ),
    .Y(\soc/cpu/_03258_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07876_  (.A(\soc/cpu/_01421_ ),
    .B(\soc/cpu/_03258_ ),
    .Y(\soc/cpu/_03259_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07877_  (.A1(\soc/cpu/pcpi_rs1 [27]),
    .A2(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03260_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_07878_  (.A1(\soc/cpu/_03227_ ),
    .A2(\soc/cpu/_03259_ ),
    .B1(\soc/cpu/_03260_ ),
    .B2(\soc/cpu/_03222_ ),
    .Y(\soc/cpu/_03261_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07879_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03257_ ),
    .B1(\soc/cpu/_03261_ ),
    .Y(\soc/cpu/_03262_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07880_  (.A(\soc/cpu/pcpi_rs1 [28]),
    .B(net47),
    .Y(\soc/cpu/_03263_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07881_  (.A1(net47),
    .A2(\soc/cpu/_03254_ ),
    .A3(\soc/cpu/_03262_ ),
    .B1(\soc/cpu/_03263_ ),
    .Y(\soc/cpu/_00698_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07882_  (.A(\soc/cpu/_02611_ ),
    .B(\soc/cpu/_02685_ ),
    .Y(\soc/cpu/_03264_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07883_  (.A1(\soc/cpu/_02684_ ),
    .A2(\soc/cpu/_03264_ ),
    .B1(\soc/cpu/_00838_ ),
    .Y(\soc/cpu/_03265_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07884_  (.A1(\soc/cpu/_02684_ ),
    .A2(\soc/cpu/_03264_ ),
    .B1(\soc/cpu/_03265_ ),
    .Y(\soc/cpu/_03266_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07885_  (.A(\soc/cpu/cpuregs_rdata1[29] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03267_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07886_  (.A(\soc/cpu/reg_pc[29] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03268_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07887_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03267_ ),
    .B1(\soc/cpu/_03268_ ),
    .Y(\soc/cpu/_03269_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07888_  (.A1(\soc/cpu/pcpi_rs1 [28]),
    .A2(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03270_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/_07889_  (.A1(\soc/cpu/_03236_ ),
    .A2(\soc/cpu/_03259_ ),
    .B1(\soc/cpu/_03270_ ),
    .B2(\soc/cpu/_03235_ ),
    .Y(\soc/cpu/_03271_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07890_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03269_ ),
    .B1(\soc/cpu/_03271_ ),
    .Y(\soc/cpu/_03272_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07891_  (.A(\soc/cpu/pcpi_rs1 [29]),
    .B(net47),
    .Y(\soc/cpu/_03273_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07892_  (.A1(net47),
    .A2(\soc/cpu/_03266_ ),
    .A3(\soc/cpu/_03272_ ),
    .B1(\soc/cpu/_03273_ ),
    .Y(\soc/cpu/_00699_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_07893_  (.A1(\soc/cpu/_02611_ ),
    .A2(\soc/cpu/_02684_ ),
    .B1(\soc/cpu/_02686_ ),
    .X(\soc/cpu/_03274_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07894_  (.A1(\soc/cpu/_02687_ ),
    .A2(\soc/cpu/_03274_ ),
    .B1(\soc/cpu/_01429_ ),
    .Y(\soc/cpu/_03275_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_07895_  (.A_N(\soc/cpu/_03275_ ),
    .B(\soc/cpu/_02688_ ),
    .Y(\soc/cpu/_03276_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07896_  (.A(\soc/cpu/cpuregs_rdata1[30] ),
    .B(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03277_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07897_  (.A(\soc/cpu/reg_pc[30] ),
    .B(\soc/cpu/_02699_ ),
    .Y(\soc/cpu/_03278_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_07898_  (.A1(\soc/cpu/is_lui_auipc_jal ),
    .A2(\soc/cpu/_03277_ ),
    .B1(\soc/cpu/_03278_ ),
    .Y(\soc/cpu/_03279_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07899_  (.A1(\soc/cpu/pcpi_rs1 [29]),
    .A2(\soc/cpu/_02603_ ),
    .B1(\soc/cpu/_02950_ ),
    .Y(\soc/cpu/_03280_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_07900_  (.A1(\soc/cpu/_03247_ ),
    .A2(\soc/cpu/_03259_ ),
    .B1(\soc/cpu/_03280_ ),
    .B2(\soc/cpu/_03246_ ),
    .Y(\soc/cpu/_03281_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07901_  (.A1(\soc/cpu/_02692_ ),
    .A2(\soc/cpu/_03279_ ),
    .B1(\soc/cpu/_03281_ ),
    .Y(\soc/cpu/_03282_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07902_  (.A(\soc/cpu/pcpi_rs1 [30]),
    .B(net47),
    .Y(\soc/cpu/_03283_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_07903_  (.A1(net47),
    .A2(\soc/cpu/_03276_ ),
    .A3(\soc/cpu/_03282_ ),
    .B1(\soc/cpu/_03283_ ),
    .Y(\soc/cpu/_00700_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07904_  (.A1(\soc/cpu/_00721_ ),
    .A2(\soc/cpu/_00825_ ),
    .B1(\soc/cpu/_00723_ ),
    .Y(\soc/cpu/_00075_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07905_  (.A1(\soc/cpu/_00721_ ),
    .A2(\soc/cpu/_00826_ ),
    .B1(\soc/cpu/_00732_ ),
    .Y(\soc/cpu/_00076_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07906_  (.A(\soc/cpu/_00718_ ),
    .B(\soc/cpu/_01110_ ),
    .Y(\soc/cpu/_03284_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07907_  (.A(\soc/cpu/_01106_ ),
    .B(\soc/cpu/_03284_ ),
    .Y(\soc/cpu/_00077_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07908_  (.A1(net65),
    .A2(\soc/cpu/_01241_ ),
    .B1(\soc/cpu/_01111_ ),
    .Y(\soc/cpu/_00078_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07909_  (.A1(\soc/cpu/_00721_ ),
    .A2(\soc/cpu/_01102_ ),
    .B1(\soc/cpu/_01096_ ),
    .Y(\soc/cpu/_00079_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07910_  (.A1(net66),
    .A2(\soc/cpu/_01088_ ),
    .B1(\soc/cpu/_01082_ ),
    .Y(\soc/cpu/_00080_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07911_  (.A1(net66),
    .A2(\soc/cpu/_01095_ ),
    .B1(\soc/cpu/_01089_ ),
    .Y(\soc/cpu/_00081_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07912_  (.A(\soc/cpu/_02351_ ),
    .B(\soc/cpu/_02354_ ),
    .Y(\soc/cpu/_03285_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07913_  (.A(\soc/cpu/prefetched_high_word ),
    .B(\soc/cpu/_03285_ ),
    .Y(\soc/cpu/_03286_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_07914_  (.A(\soc/cpu/_02351_ ),
    .Y(\soc/cpu/_03287_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_07915_  (.A(\soc/cpu/_03287_ ),
    .B(\soc/cpu/_02355_ ),
    .X(\soc/cpu/_03288_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07916_  (.A1(\soc/cpu/_03286_ ),
    .A2(\soc/cpu/_03288_ ),
    .B1(\soc/cpu/trap ),
    .C1(\soc/cpu/clear_prefetched_high_word ),
    .Y(\soc/cpu/_00099_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_07917_  (.A(\soc/cpu/irq_state[1] ),
    .B(\soc/cpu/irq_state[0] ),
    .C(\soc/cpu/_00790_ ),
    .Y(\soc/cpu/_03289_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07918_  (.A(\soc/cpu/irq_pending[20] ),
    .B(\soc/cpu/irq_pending[21] ),
    .C(\soc/cpu/irq_pending[22] ),
    .D(\soc/cpu/irq_pending[23] ),
    .Y(\soc/cpu/_03290_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_07919_  (.A(\soc/cpu/irq_pending[16] ),
    .B(\soc/cpu/irq_pending[17] ),
    .C(\soc/cpu/irq_pending[18] ),
    .D(\soc/cpu/irq_pending[19] ),
    .Y(\soc/cpu/_03291_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07920_  (.A(\soc/cpu/irq_pending[28] ),
    .B(\soc/cpu/irq_pending[29] ),
    .C(\soc/cpu/irq_pending[30] ),
    .D(\soc/cpu/irq_pending[31] ),
    .Y(\soc/cpu/_03292_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_07921_  (.A(\soc/cpu/irq_pending[24] ),
    .B(\soc/cpu/irq_pending[25] ),
    .C(\soc/cpu/irq_pending[26] ),
    .D(\soc/cpu/irq_pending[27] ),
    .Y(\soc/cpu/_03293_ ));
 sky130_fd_sc_hd__nand4_4 \soc/cpu/_07922_  (.A(\soc/cpu/_03290_ ),
    .B(\soc/cpu/_03291_ ),
    .C(\soc/cpu/_03292_ ),
    .D(\soc/cpu/_03293_ ),
    .Y(\soc/cpu/_03294_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07923_  (.A(\soc/cpu/irq_pending[4] ),
    .B(\soc/cpu/irq_pending[5] ),
    .C(\soc/cpu/irq_pending[6] ),
    .D(\soc/cpu/irq_pending[7] ),
    .Y(\soc/cpu/_03295_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07924_  (.A(\soc/cpu/irq_pending[0] ),
    .B(\soc/cpu/irq_pending[1] ),
    .C(\soc/cpu/irq_pending[2] ),
    .D(\soc/cpu/irq_pending[3] ),
    .Y(\soc/cpu/_03296_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07925_  (.A(\soc/cpu/irq_pending[12] ),
    .B(\soc/cpu/irq_pending[13] ),
    .C(\soc/cpu/irq_pending[14] ),
    .D(\soc/cpu/irq_pending[15] ),
    .Y(\soc/cpu/_03297_ ));
 sky130_fd_sc_hd__nor4_2 \soc/cpu/_07926_  (.A(\soc/cpu/irq_pending[8] ),
    .B(\soc/cpu/irq_pending[9] ),
    .C(\soc/cpu/irq_pending[10] ),
    .D(\soc/cpu/irq_pending[11] ),
    .Y(\soc/cpu/_03298_ ));
 sky130_fd_sc_hd__nand4_4 \soc/cpu/_07927_  (.A(\soc/cpu/_03295_ ),
    .B(\soc/cpu/_03296_ ),
    .C(\soc/cpu/_03297_ ),
    .D(\soc/cpu/_03298_ ),
    .Y(\soc/cpu/_03299_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_07928_  (.A(\soc/cpu/_00797_ ),
    .B(\soc/cpu/_03294_ ),
    .C(\soc/cpu/_03299_ ),
    .Y(\soc/cpu/_03300_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_07930_  (.A(\soc/cpu/_03289_ ),
    .B(\soc/cpu/_00859_ ),
    .C(\soc/cpu/_03300_ ),
    .X(\soc/cpu/_00165_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_07931_  (.A(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .Y(\soc/cpu/_03302_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_07932_  (.A(net132),
    .B(\soc/cpu/cpu_state[1] ),
    .Y(\soc/cpu/_03303_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07933_  (.A(\soc/cpu/_00991_ ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_03304_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07934_  (.A(_074_),
    .B(\soc/cpu/is_sll_srl_sra ),
    .Y(\soc/cpu/_03305_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07935_  (.A(\soc/cpu/is_lb_lh_lw_lbu_lhu ),
    .B(\soc/cpu/_00966_ ),
    .C(\soc/cpu/_03305_ ),
    .Y(\soc/cpu/_03306_ ));
 sky130_fd_sc_hd__o41ai_1 \soc/cpu/_07936_  (.A1(\soc/cpu/instr_rdcycle ),
    .A2(\soc/cpu/is_slli_srli_srai ),
    .A3(\soc/cpu/_00945_ ),
    .A4(\soc/cpu/_03306_ ),
    .B1(net807),
    .Y(\soc/cpu/_03307_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07937_  (.A(\soc/cpu/_00989_ ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_03308_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_07938_  (.A(\soc/cpu/_00934_ ),
    .B(\soc/cpu/_02600_ ),
    .C(\soc/cpu/_03307_ ),
    .D(\soc/cpu/_03308_ ),
    .Y(\soc/cpu/_03309_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07939_  (.A(\soc/cpu/_03294_ ),
    .B(\soc/cpu/_03299_ ),
    .Y(\soc/cpu/_03310_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_07940_  (.A(\soc/cpu/_00797_ ),
    .B(\soc/cpu/_03310_ ),
    .Y(\soc/cpu/_03311_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_07941_  (.A(\soc/cpu/instr_waitirq ),
    .B(\soc/cpu/_00926_ ),
    .Y(\soc/cpu/_03312_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07942_  (.A(\soc/cpu/_03311_ ),
    .B(\soc/cpu/_03312_ ),
    .Y(\soc/cpu/_03313_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07943_  (.A1(\soc/cpu/_00791_ ),
    .A2(\soc/cpu/_03313_ ),
    .B1(\soc/cpu/_00989_ ),
    .Y(\soc/cpu/_03314_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07944_  (.A(net396),
    .B(\soc/cpu/_00923_ ),
    .C(\soc/cpu/_03314_ ),
    .Y(\soc/cpu/_03315_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07945_  (.A1(\soc/cpu/is_sb_sh_sw ),
    .A2(\soc/cpu/_00957_ ),
    .B1(\soc/cpu/mem_do_prefetch ),
    .Y(\soc/cpu/_03316_ ));
 sky130_fd_sc_hd__a21boi_0 \soc/cpu/_07946_  (.A1(\soc/cpu/_00892_ ),
    .A2(\soc/cpu/_03316_ ),
    .B1_N(net955),
    .Y(\soc/cpu/_03317_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_07947_  (.A1(net799),
    .A2(\soc/cpu/cpu_state[4] ),
    .B1(\soc/cpu/_00989_ ),
    .C1(\soc/cpu/_03317_ ),
    .Y(\soc/cpu/_03318_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07948_  (.A(\soc/cpu/mem_do_rinst ),
    .B(\soc/cpu/_03309_ ),
    .Y(\soc/cpu/_03319_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07949_  (.A1(\soc/cpu/_03309_ ),
    .A2(\soc/cpu/_03315_ ),
    .A3(\soc/cpu/_03318_ ),
    .B1(\soc/cpu/_03319_ ),
    .Y(\soc/cpu/_03320_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07950_  (.A(\soc/cpu/_00964_ ),
    .B(\soc/cpu/_03320_ ),
    .Y(\soc/cpu/_03321_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_07951_  (.A1(\soc/cpu/_03302_ ),
    .A2(\soc/cpu/_01587_ ),
    .A3(\soc/cpu/_03304_ ),
    .B1(\soc/cpu/_03321_ ),
    .Y(\soc/cpu/_00179_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_07952_  (.A_N(\soc/cpu/instr_jal ),
    .B(\soc/cpu/decoder_trigger ),
    .Y(\soc/cpu/_03322_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_07953_  (.A(\soc/cpu/instr_waitirq ),
    .B(\soc/cpu/_03322_ ),
    .Y(\soc/cpu/_03323_ ));
 sky130_fd_sc_hd__o211a_1 \soc/cpu/_07954_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/instr_jalr ),
    .B1(\soc/cpu/_00796_ ),
    .C1(\soc/cpu/_03323_ ),
    .X(\soc/cpu/_03324_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07955_  (.A1(\soc/cpu/_00796_ ),
    .A2(\soc/cpu/_03323_ ),
    .B1(\soc/cpu/mem_do_prefetch ),
    .Y(\soc/cpu/_03325_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_07956_  (.A(net132),
    .B(\soc/cpu/_00963_ ),
    .C(\soc/cpu/_03324_ ),
    .D(\soc/cpu/_03325_ ),
    .Y(\soc/cpu/_00180_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_07957_  (.A1(\soc/cpu/_03302_ ),
    .A2(\soc/cpu/_00880_ ),
    .B1(\soc/cpu/_02411_ ),
    .C1(net132),
    .Y(\soc/cpu/_00579_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_07958_  (.A1(\soc/cpu/mem_do_rdata ),
    .A2(\soc/cpu/_00964_ ),
    .B1(\soc/cpu/_00851_ ),
    .X(\soc/cpu/_00582_ ));
 sky130_fd_sc_hd__inv_2 \soc/cpu/_07959_  (.A(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03326_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_07960_  (.A(\soc/cpu/_03326_ ),
    .B(\soc/cpu/_00989_ ),
    .Y(\soc/cpu/_03327_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_07961_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03327_ ),
    .Y(\soc/cpu/_03328_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_07963_  (.A(_074_),
    .B(\soc/cpu/_00839_ ),
    .Y(\soc/cpu/_03330_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_07964_  (.A(net778),
    .B(\soc/cpu/_00843_ ),
    .C(\soc/cpu/_03330_ ),
    .Y(\soc/cpu/_03331_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_07965_  (.A1(\soc/cpu/mem_do_wdata ),
    .A2(\soc/cpu/_00964_ ),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/_03331_ ),
    .X(\soc/cpu/_00583_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07966_  (.A1(\soc/cpu/mem_la_secondword ),
    .A2(\soc/cpu/_03287_ ),
    .B1(\soc/cpu/_02373_ ),
    .Y(\soc/cpu/_03332_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07967_  (.A(\soc/cpu/_02362_ ),
    .B(\soc/cpu/_03332_ ),
    .Y(\soc/cpu/_00100_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07968_  (.A1(\soc/cpu/_02386_ ),
    .A2(\soc/cpu/_02528_ ),
    .B1(\soc/cpu/_01279_ ),
    .Y(\soc/cpu/_03333_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07969_  (.A1(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .A2(\soc/cpu/_01588_ ),
    .B1(_074_),
    .Y(\soc/cpu/_03334_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07970_  (.A1(\soc/cpu/_01588_ ),
    .A2(\soc/cpu/_03333_ ),
    .B1(\soc/cpu/_03334_ ),
    .Y(\soc/cpu/_00108_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07971_  (.A(\soc/cpu/mem_rdata_q[0] ),
    .B(\soc/cpu/mem_rdata_q[1] ),
    .C(\soc/cpu/mem_rdata_q[2] ),
    .Y(\soc/cpu/_03335_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_07972_  (.A(\soc/cpu/_02430_ ),
    .B(\soc/cpu/_02516_ ),
    .C(\soc/cpu/_03335_ ),
    .X(\soc/cpu/_03336_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07973_  (.A1(\soc/cpu/instr_fence ),
    .A2(\soc/cpu/_02411_ ),
    .B1(_074_),
    .Y(\soc/cpu/_03337_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07974_  (.A1(\soc/cpu/_02411_ ),
    .A2(\soc/cpu/_03336_ ),
    .B1(\soc/cpu/_03337_ ),
    .Y(\soc/cpu/_00133_ ));
 sky130_fd_sc_hd__and3b_1 \soc/cpu/_07977_  (.A_N(\soc/cpu/mem_rdata_q[12] ),
    .B(net951),
    .C(net950),
    .X(\soc/cpu/_03340_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07978_  (.A(\soc/cpu/is_alu_reg_reg ),
    .B(\soc/cpu/_02411_ ),
    .Y(\soc/cpu/_03341_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/cpu/_07979_  (.A(\soc/cpu/_02419_ ),
    .SLEEP(\soc/cpu/_03341_ ),
    .X(\soc/cpu/_03342_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_07980_  (.A1(\soc/cpu/instr_or ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03340_ ),
    .B2(\soc/cpu/_03342_ ),
    .Y(\soc/cpu/_03343_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07981_  (.A(net132),
    .B(\soc/cpu/_03343_ ),
    .Y(\soc/cpu/_00136_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_07982_  (.A1(\soc/cpu/instr_srl ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02424_ ),
    .B2(\soc/cpu/_03342_ ),
    .Y(\soc/cpu/_03344_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07983_  (.A(net132),
    .B(\soc/cpu/_03344_ ),
    .Y(\soc/cpu/_00137_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_07985_  (.A1(\soc/cpu/instr_xor ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02523_ ),
    .B2(\soc/cpu/_03342_ ),
    .Y(\soc/cpu/_03346_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07986_  (.A(net132),
    .B(\soc/cpu/_03346_ ),
    .Y(\soc/cpu/_00138_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_07987_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(\soc/cpu/mem_rdata_q[13] ),
    .Y(\soc/cpu/_03347_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07988_  (.A(\soc/cpu/mem_rdata_q[14] ),
    .B(\soc/cpu/_03347_ ),
    .Y(\soc/cpu/_03348_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_07989_  (.A1(\soc/cpu/instr_sltu ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03342_ ),
    .B2(\soc/cpu/_03348_ ),
    .Y(\soc/cpu/_03349_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07990_  (.A(net132),
    .B(\soc/cpu/_03349_ ),
    .Y(\soc/cpu/_00139_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/cpu/_07991_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(net950),
    .C_N(net951),
    .Y(\soc/cpu/_03350_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_07992_  (.A1(\soc/cpu/instr_slt ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03350_ ),
    .B2(\soc/cpu/_03342_ ),
    .Y(\soc/cpu/_03351_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07993_  (.A(net132),
    .B(\soc/cpu/_03351_ ),
    .Y(\soc/cpu/_00140_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_07994_  (.A1(\soc/cpu/instr_sll ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02509_ ),
    .B2(\soc/cpu/_03342_ ),
    .Y(\soc/cpu/_03352_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_07995_  (.A(net132),
    .B(\soc/cpu/_03352_ ),
    .Y(\soc/cpu/_00141_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_07996_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(net951),
    .C(net950),
    .Y(\soc/cpu/_03353_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_07997_  (.A(net850),
    .B(\soc/cpu/_02423_ ),
    .C(\soc/cpu/_03353_ ),
    .Y(\soc/cpu/_03354_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_07998_  (.A1(\soc/cpu/instr_sub ),
    .A2(\soc/cpu/_02411_ ),
    .B1(_074_),
    .Y(\soc/cpu/_03355_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_07999_  (.A1(\soc/cpu/_02411_ ),
    .A2(\soc/cpu/_03354_ ),
    .B1(\soc/cpu/_03355_ ),
    .Y(\soc/cpu/_00142_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08000_  (.A1(\soc/cpu/instr_add ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03353_ ),
    .B2(\soc/cpu/_03342_ ),
    .Y(\soc/cpu/_03356_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08001_  (.A(net132),
    .B(\soc/cpu/_03356_ ),
    .Y(\soc/cpu/_00143_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08002_  (.A(\soc/cpu/mem_rdata_q[12] ),
    .B(net951),
    .C(net950),
    .X(\soc/cpu/_03357_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08003_  (.A1(\soc/cpu/instr_andi ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_03357_ ),
    .Y(\soc/cpu/_03358_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08004_  (.A(net132),
    .B(\soc/cpu/_03358_ ),
    .Y(\soc/cpu/_00147_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08005_  (.A1(\soc/cpu/instr_ori ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_03340_ ),
    .Y(\soc/cpu/_03359_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08006_  (.A(net132),
    .B(\soc/cpu/_03359_ ),
    .Y(\soc/cpu/_00148_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08007_  (.A1(\soc/cpu/instr_xori ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_02523_ ),
    .Y(\soc/cpu/_03360_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08008_  (.A(net132),
    .B(\soc/cpu/_03360_ ),
    .Y(\soc/cpu/_00149_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08010_  (.A1(\soc/cpu/instr_sltiu ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_03348_ ),
    .Y(\soc/cpu/_03362_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08011_  (.A(net132),
    .B(\soc/cpu/_03362_ ),
    .Y(\soc/cpu/_00150_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08012_  (.A1(\soc/cpu/instr_slti ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_03350_ ),
    .Y(\soc/cpu/_03363_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08013_  (.A(net132),
    .B(\soc/cpu/_03363_ ),
    .Y(\soc/cpu/_00151_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08014_  (.A1(\soc/cpu/instr_addi ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02412_ ),
    .B2(\soc/cpu/_03353_ ),
    .Y(\soc/cpu/_03364_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08015_  (.A(net132),
    .B(\soc/cpu/_03364_ ),
    .Y(\soc/cpu/_00152_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_08016_  (.A(\soc/cpu/_03302_ ),
    .B(\soc/cpu/_02408_ ),
    .Y(\soc/cpu/_03365_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08017_  (.A1(\soc/cpu/instr_bltu ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03340_ ),
    .B2(\soc/cpu/_03365_ ),
    .Y(\soc/cpu/_03366_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08018_  (.A(net132),
    .B(\soc/cpu/_03366_ ),
    .Y(\soc/cpu/_00159_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08019_  (.A1(\soc/cpu/instr_bge ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02424_ ),
    .B2(\soc/cpu/_03365_ ),
    .Y(\soc/cpu/_03367_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08020_  (.A(net132),
    .B(\soc/cpu/_03367_ ),
    .Y(\soc/cpu/_00160_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08021_  (.A1(\soc/cpu/instr_blt ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02523_ ),
    .B2(\soc/cpu/_03365_ ),
    .Y(\soc/cpu/_03368_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08022_  (.A(net132),
    .B(\soc/cpu/_03368_ ),
    .Y(\soc/cpu/_00161_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08023_  (.A1(\soc/cpu/instr_bne ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_02509_ ),
    .B2(\soc/cpu/_03365_ ),
    .Y(\soc/cpu/_03369_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08024_  (.A(net132),
    .B(\soc/cpu/_03369_ ),
    .Y(\soc/cpu/_00162_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_08025_  (.A(\soc/cpu/_00839_ ),
    .B(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03370_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08026_  (.A1(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .A2(\soc/cpu/cpu_state[3] ),
    .B1(\soc/cpu/_03370_ ),
    .Y(\soc/cpu/_03371_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08027_  (.A(\soc/cpu/cpuregs_waddr[0] ),
    .B(\soc/cpu/_03371_ ),
    .Y(\soc/cpu/_03372_ ));
 sky130_fd_sc_hd__o311ai_1 \soc/cpu/_08028_  (.A1(\soc/cpu/irq_state[1] ),
    .A2(\soc/cpu/decoded_rd[0] ),
    .A3(\soc/cpu/_00790_ ),
    .B1(\soc/cpu/_03370_ ),
    .C1(\soc/cpu/_02143_ ),
    .Y(\soc/cpu/_03373_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08030_  (.A1(\soc/cpu/_03372_ ),
    .A2(\soc/cpu/_03373_ ),
    .B1(net132),
    .Y(\soc/cpu/_00167_ ));
 sky130_fd_sc_hd__o311ai_1 \soc/cpu/_08032_  (.A1(\soc/cpu/irq_state[1] ),
    .A2(\soc/cpu/decoded_rd[1] ),
    .A3(\soc/cpu/_00790_ ),
    .B1(\soc/cpu/_03370_ ),
    .C1(\soc/cpu/_02143_ ),
    .Y(\soc/cpu/_03376_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08033_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/_03371_ ),
    .Y(\soc/cpu/_03377_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08034_  (.A(_074_),
    .B(\soc/cpu/_03376_ ),
    .C(\soc/cpu/_03377_ ),
    .Y(\soc/cpu/_00168_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08035_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/decoded_rd[2] ),
    .B1(\soc/cpu/_03370_ ),
    .Y(\soc/cpu/_03378_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08036_  (.A1(\soc/cpu/_02143_ ),
    .A2(\soc/cpu/_00791_ ),
    .B1(\soc/cpu/_03378_ ),
    .Y(\soc/cpu/_03379_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08037_  (.A1(\soc/cpu/cpuregs_waddr[2] ),
    .A2(\soc/cpu/_03371_ ),
    .B1(\soc/cpu/_03379_ ),
    .Y(\soc/cpu/_03380_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08038_  (.A(net132),
    .B(\soc/cpu/_03380_ ),
    .Y(\soc/cpu/_00169_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08039_  (.A(_074_),
    .B(\soc/cpu/_03289_ ),
    .Y(\soc/cpu/_03381_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08040_  (.A(\soc/cpu/decoded_rd[3] ),
    .B(\soc/cpu/_03370_ ),
    .Y(\soc/cpu/_03382_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08041_  (.A(_074_),
    .B(\soc/cpu/cpuregs_waddr[3] ),
    .C(\soc/cpu/_03371_ ),
    .Y(\soc/cpu/_03383_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08042_  (.A1(\soc/cpu/_03381_ ),
    .A2(\soc/cpu/_03382_ ),
    .B1(\soc/cpu/_03383_ ),
    .Y(\soc/cpu/_00170_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08043_  (.A(net898),
    .B(\soc/cpu/_03370_ ),
    .Y(\soc/cpu/_03384_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08044_  (.A(_074_),
    .B(\soc/cpu/cpuregs_waddr[4] ),
    .C(\soc/cpu/_03371_ ),
    .Y(\soc/cpu/_03385_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08045_  (.A1(\soc/cpu/_03381_ ),
    .A2(\soc/cpu/_03384_ ),
    .B1(\soc/cpu/_03385_ ),
    .Y(\soc/cpu/_00171_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08046_  (.A(\soc/cpu/cpu_state[6] ),
    .B(net800),
    .Y(\soc/cpu/_03386_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_08047_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/cpu_state[6] ),
    .B1(\soc/cpu/_03386_ ),
    .B2(\soc/cpu/mem_do_rdata ),
    .Y(\soc/cpu/_03387_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08048_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/instr_lb ),
    .Y(\soc/cpu/_03388_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08049_  (.A(\soc/cpu/latched_is_lb ),
    .B(\soc/cpu/_03387_ ),
    .Y(\soc/cpu/_03389_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_08050_  (.A1(\soc/cpu/_03387_ ),
    .A2(\soc/cpu/_03388_ ),
    .B1(\soc/cpu/_03389_ ),
    .C1(net132),
    .Y(\soc/cpu/_00172_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08051_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/instr_lh ),
    .Y(\soc/cpu/_03390_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08052_  (.A(\soc/cpu/latched_is_lh ),
    .B(\soc/cpu/_03387_ ),
    .Y(\soc/cpu/_03391_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_08053_  (.A1(\soc/cpu/_03387_ ),
    .A2(\soc/cpu/_03390_ ),
    .B1(\soc/cpu/_03391_ ),
    .C1(net132),
    .Y(\soc/cpu/_00173_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08054_  (.A1(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .A2(\soc/cpu/_01587_ ),
    .B1(\soc/cpu/_00940_ ),
    .Y(\soc/cpu/_03392_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08055_  (.A1(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .A2(\soc/cpu/instr_jalr ),
    .B1(\soc/cpu/_03392_ ),
    .Y(\soc/cpu/_03393_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08057_  (.A(net413),
    .B(\soc/cpu/cpu_state[1] ),
    .C(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03395_ ));
 sky130_fd_sc_hd__a311oi_1 \soc/cpu/_08058_  (.A1(\soc/cpu/_00940_ ),
    .A2(\soc/cpu/_03289_ ),
    .A3(\soc/cpu/_03312_ ),
    .B1(\soc/cpu/_03395_ ),
    .C1(net413),
    .Y(\soc/cpu/_03396_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_08059_  (.A(net413),
    .SLEEP(\soc/cpu/instr_retirq ),
    .X(\soc/cpu/_03397_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08060_  (.A1(\soc/cpu/_03395_ ),
    .A2(\soc/cpu/_03397_ ),
    .B1(\soc/cpu/_02108_ ),
    .Y(\soc/cpu/_03398_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08061_  (.A(_074_),
    .B(\soc/cpu/_03398_ ),
    .Y(\soc/cpu/_03399_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08062_  (.A1(\soc/cpu/_03393_ ),
    .A2(\soc/cpu/_03396_ ),
    .B1(\soc/cpu/_03399_ ),
    .Y(\soc/cpu/_00175_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_08065_  (.A1(net807),
    .A2(\soc/cpu/_00946_ ),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/_00839_ ),
    .Y(\soc/cpu/_03402_ ));
 sky130_fd_sc_hd__clkinv_4 \soc/cpu/_08066_  (.A(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_03403_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08067_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_00791_ ),
    .C(\soc/cpu/_03403_ ),
    .Y(\soc/cpu/_03404_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_08068_  (.A1(\soc/cpu/_03327_ ),
    .A2(\soc/cpu/_03392_ ),
    .A3(\soc/cpu/_03404_ ),
    .B1(\soc/cpu/_03402_ ),
    .Y(\soc/cpu/_03405_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_08069_  (.A1(\soc/cpu/_00985_ ),
    .A2(\soc/cpu/_03402_ ),
    .B1(\soc/cpu/_03405_ ),
    .C1(_074_),
    .Y(\soc/cpu/_00176_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/_08071_  (.A(\soc/cpu/irq_state[1] ),
    .B(\soc/cpu/cpu_state[1] ),
    .Y(\soc/cpu/_03407_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08072_  (.A(\soc/cpu/irq_state[0] ),
    .B(net819),
    .Y(\soc/cpu/_03408_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08073_  (.A(_074_),
    .B(\soc/cpu/_03407_ ),
    .C(\soc/cpu/_03408_ ),
    .Y(\soc/cpu/_03409_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08074_  (.A1(\soc/cpu/_02143_ ),
    .A2(\soc/cpu/_00953_ ),
    .B1(\soc/cpu/_03409_ ),
    .Y(\soc/cpu/_00177_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08076_  (.A(_074_),
    .B(\soc/cpu/_03407_ ),
    .Y(\soc/cpu/_03411_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08077_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(net819),
    .B1(\soc/cpu/irq_state[1] ),
    .Y(\soc/cpu/_03412_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08078_  (.A(\soc/cpu/_03411_ ),
    .B(\soc/cpu/_03412_ ),
    .Y(\soc/cpu/_00178_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_16 \soc/cpu/_08080_  (.A(net160),
    .SLEEP(\soc/cpu/_00873_ ),
    .X(\soc/cpu/_03414_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08082_  (.A1(\soc/cpu/count_instr[0] ),
    .A2(\soc/cpu/instr_rdinstr ),
    .B1(\soc/cpu/instr_rdcycleh ),
    .B2(\soc/cpu/count_cycle[32] ),
    .C1(\soc/cpu/count_instr[32] ),
    .C2(\soc/cpu/instr_rdinstrh ),
    .Y(\soc/cpu/_03416_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08083_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03416_ ),
    .Y(\soc/cpu/_03417_ ));
 sky130_fd_sc_hd__a221o_2 \soc/cpu/_08085_  (.A1(\soc/cpu/irq_mask[0] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[0] ),
    .C1(\soc/cpu/_00872_ ),
    .X(\soc/cpu/_03419_ ));
 sky130_fd_sc_hd__o2111ai_4 \soc/cpu/_08086_  (.A1(\soc/cpu/count_cycle[0] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03417_ ),
    .C1(\soc/cpu/_03419_ ),
    .D1(net413),
    .Y(\soc/cpu/_03420_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08088_  (.A1(\soc/cpu/reg_next_pc[0] ),
    .A2(\soc/cpu/decoded_imm[0] ),
    .B1(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03422_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08089_  (.A1(\soc/cpu/reg_next_pc[0] ),
    .A2(\soc/cpu/decoded_imm[0] ),
    .B1(\soc/cpu/_03422_ ),
    .Y(\soc/cpu/_03423_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08090_  (.A1(\soc/cpu/pcpi_rs1 [0]),
    .A2(\soc/cpu/cpu_state[4] ),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[0] ),
    .C1(\soc/cpu/_03423_ ),
    .Y(\soc/cpu/_03424_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/_08091_  (.A0(\soc/mem_rdata[8] ),
    .A1(\soc/mem_rdata[24] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .Y(\soc/cpu/_03425_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08092_  (.A(\soc/cpu/pcpi_rs1 [0]),
    .B(\soc/cpu/mem_wordsize[1] ),
    .Y(\soc/cpu/_03426_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08093_  (.A(\soc/cpu/mem_wordsize[1] ),
    .B(\soc/cpu/_02285_ ),
    .Y(\soc/cpu/_03427_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_08094_  (.A(\soc/cpu/_02282_ ),
    .B(\soc/cpu/_03427_ ),
    .Y(\soc/cpu/_03428_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08095_  (.A1(\soc/mem_rdata[0] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03428_ ),
    .B2(\soc/mem_rdata[16] ),
    .Y(\soc/cpu/_03429_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08096_  (.A1(\soc/cpu/_03425_ ),
    .A2(\soc/cpu/_03426_ ),
    .B1(\soc/cpu/_03429_ ),
    .Y(\soc/cpu/_03430_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08097_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/_03430_ ),
    .Y(\soc/cpu/_03431_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08099_  (.A1(\soc/cpu/_03420_ ),
    .A2(\soc/cpu/_03424_ ),
    .A3(\soc/cpu/_03431_ ),
    .B1(net132),
    .Y(\soc/cpu/_00181_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08101_  (.A(\soc/cpu/decoded_imm[1] ),
    .B(\soc/cpu/reg_pc[1] ),
    .Y(\soc/cpu/_03434_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08102_  (.A(\soc/cpu/decoded_imm[1] ),
    .B(\soc/cpu/reg_pc[1] ),
    .X(\soc/cpu/_03435_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08103_  (.A(\soc/cpu/reg_next_pc[0] ),
    .B(\soc/cpu/decoded_imm[0] ),
    .Y(\soc/cpu/_03436_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08104_  (.A1(\soc/cpu/_03434_ ),
    .A2(\soc/cpu/_03435_ ),
    .B1(\soc/cpu/_03436_ ),
    .Y(\soc/cpu/_03437_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_08105_  (.A(\soc/cpu/_03436_ ),
    .B(\soc/cpu/_03434_ ),
    .C(\soc/cpu/_03435_ ),
    .X(\soc/cpu/_03438_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_08106_  (.A0(\soc/mem_rdata[9] ),
    .A1(\soc/mem_rdata[25] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .Y(\soc/cpu/_03439_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08107_  (.A(\soc/cpu/_03426_ ),
    .B(\soc/cpu/_03439_ ),
    .Y(\soc/cpu/_03440_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08108_  (.A1(\soc/mem_rdata[1] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03428_ ),
    .B2(\soc/mem_rdata[17] ),
    .C1(\soc/cpu/_03440_ ),
    .Y(\soc/cpu/_03441_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08109_  (.A1(\soc/cpu/pcpi_rs1 [1]),
    .A2(\soc/cpu/cpu_state[4] ),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[1] ),
    .Y(\soc/cpu/_03442_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08110_  (.A1(\soc/cpu/_03326_ ),
    .A2(\soc/cpu/_03441_ ),
    .B1(\soc/cpu/_03442_ ),
    .Y(\soc/cpu/_03443_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08111_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03437_ ),
    .A3(\soc/cpu/_03438_ ),
    .B1(\soc/cpu/_03443_ ),
    .Y(\soc/cpu/_03444_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_08113_  (.A_N(\soc/cpu/_00873_ ),
    .B(net160),
    .Y(\soc/cpu/_03446_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08115_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[33] ),
    .B1(\soc/cpu/count_instr[1] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[33] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03448_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08116_  (.A(\soc/cpu/_02935_ ),
    .Y(\soc/cpu/_03449_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08117_  (.A1(\soc/cpu/irq_mask[1] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[1] ),
    .C1(\soc/cpu/_03449_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03450_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08118_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03448_ ),
    .B1(\soc/cpu/_03450_ ),
    .Y(\soc/cpu/_03451_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08119_  (.A1(\soc/cpu/count_cycle[1] ),
    .A2(\soc/cpu/_00874_ ),
    .B1(\soc/cpu/_03451_ ),
    .Y(\soc/cpu/_03452_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_08120_  (.A1(net132),
    .A2(\soc/cpu/_03444_ ),
    .B1(\soc/cpu/_03452_ ),
    .B2(\soc/cpu/_00894_ ),
    .Y(\soc/cpu/_00182_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08121_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[34] ),
    .B1(\soc/cpu/count_instr[2] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[34] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03453_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08122_  (.A(\soc/cpu/count_cycle[2] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03454_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08123_  (.A(\soc/cpu/_02945_ ),
    .Y(\soc/cpu/_03455_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08124_  (.A1(\soc/cpu/irq_mask[2] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[2] ),
    .C1(\soc/cpu/_03455_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03456_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_08125_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03453_ ),
    .B1(\soc/cpu/_03454_ ),
    .C1(\soc/cpu/_03456_ ),
    .Y(\soc/cpu/_03457_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_08126_  (.A(net413),
    .B(\soc/cpu/_03457_ ),
    .Y(\soc/cpu/_03458_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08127_  (.A(\soc/mem_rdata[2] ),
    .B(\soc/cpu/mem_la_wstrb [0]),
    .Y(\soc/cpu/_03459_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_08128_  (.A0(\soc/mem_rdata[10] ),
    .A1(\soc/mem_rdata[26] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .X(\soc/cpu/_03460_ ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_08129_  (.A(\soc/cpu/pcpi_rs1 [0]),
    .B(\soc/cpu/mem_wordsize[1] ),
    .X(\soc/cpu/_03461_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08130_  (.A1(\soc/mem_rdata[18] ),
    .A2(\soc/cpu/_03428_ ),
    .B1(\soc/cpu/_03460_ ),
    .B2(\soc/cpu/_03461_ ),
    .Y(\soc/cpu/_03462_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08131_  (.A(\soc/cpu/_03459_ ),
    .B(\soc/cpu/_03462_ ),
    .Y(\soc/cpu/_03463_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08132_  (.A(\soc/cpu/cpu_state[6] ),
    .B(\soc/cpu/_03463_ ),
    .Y(\soc/cpu/_03464_ ));
 sky130_fd_sc_hd__o21ba_1 \soc/cpu/_08133_  (.A1(\soc/cpu/_03436_ ),
    .A2(\soc/cpu/_03434_ ),
    .B1_N(\soc/cpu/_03435_ ),
    .X(\soc/cpu/_03465_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08134_  (.A(\soc/cpu/decoded_imm[2] ),
    .B(\soc/cpu/reg_pc[2] ),
    .Y(\soc/cpu/_03466_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_08135_  (.A(\soc/cpu/_03465_ ),
    .B(\soc/cpu/_03466_ ),
    .X(\soc/cpu/_03467_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08136_  (.A1(\soc/cpu/irq_pending[2] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03467_ ),
    .B2(\soc/cpu/cpu_state[3] ),
    .C1(\soc/cpu/cpu_state[4] ),
    .C2(\soc/cpu/pcpi_rs1 [2]),
    .Y(\soc/cpu/_03468_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08137_  (.A1(\soc/cpu/_03458_ ),
    .A2(\soc/cpu/_03464_ ),
    .A3(\soc/cpu/_03468_ ),
    .B1(net132),
    .Y(\soc/cpu/_00183_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08138_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[3] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03469_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08139_  (.A1(\soc/cpu/irq_mask[3] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[3] ),
    .C1(net160),
    .Y(\soc/cpu/_03470_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08140_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[35] ),
    .B1(\soc/cpu/count_instr[3] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[35] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03471_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08141_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03471_ ),
    .Y(\soc/cpu/_03472_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08142_  (.A1(\soc/cpu/count_cycle[3] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03472_ ),
    .Y(\soc/cpu/_03473_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08143_  (.A1(\soc/cpu/_03469_ ),
    .A2(\soc/cpu/_03470_ ),
    .B1(\soc/cpu/_03473_ ),
    .Y(\soc/cpu/_03474_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_08144_  (.A0(\soc/mem_rdata[11] ),
    .A1(\soc/mem_rdata[27] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .X(\soc/cpu/_03475_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08145_  (.A1(\soc/mem_rdata[3] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03461_ ),
    .B2(\soc/cpu/_03475_ ),
    .C1(\soc/cpu/_03428_ ),
    .C2(\soc/mem_rdata[19] ),
    .Y(\soc/cpu/_03476_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08147_  (.A(\soc/cpu/decoded_imm[2] ),
    .B(\soc/cpu/reg_pc[2] ),
    .Y(\soc/cpu/_03478_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08148_  (.A1(\soc/cpu/_03465_ ),
    .A2(\soc/cpu/_03466_ ),
    .B1(\soc/cpu/_03478_ ),
    .Y(\soc/cpu/_03479_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08149_  (.A(\soc/cpu/decoded_imm[3] ),
    .B(\soc/cpu/reg_pc[3] ),
    .Y(\soc/cpu/_03480_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08150_  (.A(\soc/cpu/decoded_imm[3] ),
    .B(\soc/cpu/reg_pc[3] ),
    .Y(\soc/cpu/_03481_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_08151_  (.A_N(\soc/cpu/_03480_ ),
    .B(\soc/cpu/_03481_ ),
    .Y(\soc/cpu/_03482_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08152_  (.A(\soc/cpu/_03479_ ),
    .B(\soc/cpu/_03482_ ),
    .Y(\soc/cpu/_03483_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08153_  (.A1(\soc/cpu/irq_pending[3] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03483_ ),
    .B2(\soc/cpu/cpu_state[3] ),
    .C1(\soc/cpu/cpu_state[4] ),
    .C2(\soc/cpu/pcpi_rs1 [3]),
    .Y(\soc/cpu/_03484_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08154_  (.A1(\soc/cpu/_03326_ ),
    .A2(\soc/cpu/_03476_ ),
    .B1(\soc/cpu/_03484_ ),
    .Y(\soc/cpu/_03485_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08155_  (.A1(\soc/cpu/cpu_state[2] ),
    .A2(\soc/cpu/_03474_ ),
    .B1(\soc/cpu/_03485_ ),
    .Y(\soc/cpu/_03486_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08156_  (.A(net132),
    .B(\soc/cpu/_03486_ ),
    .Y(\soc/cpu/_00184_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_08157_  (.A(\soc/cpu/decoded_imm[4] ),
    .B(\soc/cpu/reg_pc[4] ),
    .Y(\soc/cpu/_03487_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08158_  (.A1(\soc/cpu/decoded_imm[3] ),
    .A2(\soc/cpu/reg_pc[3] ),
    .B1(\soc/cpu/_03479_ ),
    .Y(\soc/cpu/_03488_ ));
 sky130_fd_sc_hd__o211a_1 \soc/cpu/_08159_  (.A1(\soc/cpu/_03465_ ),
    .A2(\soc/cpu/_03466_ ),
    .B1(\soc/cpu/_03481_ ),
    .C1(\soc/cpu/_03478_ ),
    .X(\soc/cpu/_03489_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_08160_  (.A1(\soc/cpu/_03480_ ),
    .A2(\soc/cpu/_03487_ ),
    .A3(\soc/cpu/_03489_ ),
    .B1(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03490_ ));
 sky130_fd_sc_hd__a31o_1 \soc/cpu/_08161_  (.A1(\soc/cpu/_03481_ ),
    .A2(\soc/cpu/_03487_ ),
    .A3(\soc/cpu/_03488_ ),
    .B1(\soc/cpu/_03490_ ),
    .X(\soc/cpu/_03491_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08162_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [4]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[4] ),
    .Y(\soc/cpu/_03492_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08166_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[36] ),
    .B1(\soc/cpu/count_instr[4] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[36] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03496_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08167_  (.A(\soc/cpu/count_cycle[4] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03497_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08170_  (.A(\soc/cpu/_02980_ ),
    .Y(\soc/cpu/_03500_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08172_  (.A1(\soc/cpu/irq_mask[4] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[4] ),
    .C1(\soc/cpu/_03500_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03502_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08173_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03496_ ),
    .B1(\soc/cpu/_03497_ ),
    .C1(\soc/cpu/_03502_ ),
    .Y(\soc/cpu/_03503_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_08174_  (.A0(\soc/mem_rdata[12] ),
    .A1(\soc/mem_rdata[28] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .X(\soc/cpu/_03504_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08175_  (.A1(\soc/mem_rdata[4] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03461_ ),
    .B2(\soc/cpu/_03504_ ),
    .C1(\soc/cpu/_03428_ ),
    .C2(\soc/mem_rdata[20] ),
    .Y(\soc/cpu/_03505_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08176_  (.A(\soc/cpu/_03326_ ),
    .B(\soc/cpu/_03505_ ),
    .Y(\soc/cpu/_03506_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08177_  (.A1(\soc/cpu/cpu_state[2] ),
    .A2(\soc/cpu/_03503_ ),
    .B1(\soc/cpu/_03506_ ),
    .Y(\soc/cpu/_03507_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_08178_  (.A1(\soc/cpu/_03491_ ),
    .A2(\soc/cpu/_03492_ ),
    .A3(\soc/cpu/_03507_ ),
    .B1(net132),
    .Y(\soc/cpu/_00185_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08179_  (.A(\soc/cpu/decoded_imm[4] ),
    .B(\soc/cpu/reg_pc[4] ),
    .Y(\soc/cpu/_03508_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_08180_  (.A1(\soc/cpu/_03480_ ),
    .A2(\soc/cpu/_03487_ ),
    .A3(\soc/cpu/_03489_ ),
    .B1(\soc/cpu/_03508_ ),
    .Y(\soc/cpu/_03509_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_08181_  (.A(\soc/cpu/decoded_imm[5] ),
    .B(\soc/cpu/reg_pc[5] ),
    .X(\soc/cpu/_03510_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08182_  (.A(\soc/cpu/decoded_imm[5] ),
    .B(\soc/cpu/reg_pc[5] ),
    .Y(\soc/cpu/_03511_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08183_  (.A(\soc/cpu/_03510_ ),
    .B(\soc/cpu/_03511_ ),
    .Y(\soc/cpu/_03512_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08184_  (.A(\soc/cpu/_03509_ ),
    .B(\soc/cpu/_03512_ ),
    .Y(\soc/cpu/_03513_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_08185_  (.A0(\soc/mem_rdata[13] ),
    .A1(\soc/mem_rdata[29] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .X(\soc/cpu/_03514_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08186_  (.A1(\soc/mem_rdata[5] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03461_ ),
    .B2(\soc/cpu/_03514_ ),
    .C1(\soc/cpu/_03428_ ),
    .C2(\soc/mem_rdata[21] ),
    .Y(\soc/cpu/_03515_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08189_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[5] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03518_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08192_  (.A1(\soc/cpu/irq_mask[5] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[5] ),
    .C1(net160),
    .Y(\soc/cpu/_03521_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08198_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[37] ),
    .B1(\soc/cpu/count_instr[5] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[37] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03527_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08199_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03527_ ),
    .Y(\soc/cpu/_03528_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08200_  (.A1(\soc/cpu/count_cycle[5] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03528_ ),
    .Y(\soc/cpu/_03529_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08201_  (.A1(\soc/cpu/_03518_ ),
    .A2(\soc/cpu/_03521_ ),
    .B1(\soc/cpu/_03529_ ),
    .Y(\soc/cpu/_03530_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08202_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [5]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[5] ),
    .C1(net413),
    .C2(\soc/cpu/_03530_ ),
    .Y(\soc/cpu/_03531_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08203_  (.A1(\soc/cpu/_03326_ ),
    .A2(\soc/cpu/_03515_ ),
    .B1(\soc/cpu/_03531_ ),
    .Y(\soc/cpu/_03532_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08204_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03513_ ),
    .B1(\soc/cpu/_03532_ ),
    .Y(\soc/cpu/_03533_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08205_  (.A(net132),
    .B(\soc/cpu/_03533_ ),
    .Y(\soc/cpu/_00186_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08207_  (.A1(\soc/cpu/_03509_ ),
    .A2(\soc/cpu/_03510_ ),
    .B1_N(\soc/cpu/_03511_ ),
    .Y(\soc/cpu/_03535_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08208_  (.A(\soc/cpu/decoded_imm[6] ),
    .B(\soc/cpu/reg_pc[6] ),
    .Y(\soc/cpu/_03536_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08209_  (.A(\soc/cpu/_03535_ ),
    .B(\soc/cpu/_03536_ ),
    .Y(\soc/cpu/_03537_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_08210_  (.A(\soc/cpu/_03535_ ),
    .B(\soc/cpu/_03536_ ),
    .X(\soc/cpu/_03538_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08211_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03537_ ),
    .C(\soc/cpu/_03538_ ),
    .Y(\soc/cpu/_03539_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08212_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [6]),
    .B1(\soc/cpu/_03328_ ),
    .B2(net960),
    .Y(\soc/cpu/_03540_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08213_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[38] ),
    .B1(\soc/cpu/count_instr[6] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[38] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03541_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08214_  (.A(\soc/cpu/count_cycle[6] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03542_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08215_  (.A(\soc/cpu/_03008_ ),
    .Y(\soc/cpu/_03543_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08216_  (.A1(\soc/cpu/irq_mask[6] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[6] ),
    .C1(\soc/cpu/_03543_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03544_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08217_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03541_ ),
    .B1(\soc/cpu/_03542_ ),
    .C1(\soc/cpu/_03544_ ),
    .Y(\soc/cpu/_03545_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/_08218_  (.A0(\soc/mem_rdata[14] ),
    .A1(\soc/mem_rdata[30] ),
    .S(\soc/cpu/pcpi_rs1 [1]),
    .X(\soc/cpu/_03546_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08219_  (.A1(\soc/mem_rdata[6] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03461_ ),
    .B2(\soc/cpu/_03546_ ),
    .C1(\soc/cpu/_03428_ ),
    .C2(\soc/mem_rdata[22] ),
    .Y(\soc/cpu/_03547_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08220_  (.A(\soc/cpu/_03326_ ),
    .B(\soc/cpu/_03547_ ),
    .Y(\soc/cpu/_03548_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08221_  (.A1(net801),
    .A2(\soc/cpu/_03545_ ),
    .B1(\soc/cpu/_03548_ ),
    .Y(\soc/cpu/_03549_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08222_  (.A1(\soc/cpu/_03539_ ),
    .A2(net961),
    .A3(\soc/cpu/_03549_ ),
    .B1(net131),
    .Y(\soc/cpu/_00187_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08223_  (.A(\soc/cpu/decoded_imm[6] ),
    .B(\soc/cpu/reg_pc[6] ),
    .Y(\soc/cpu/_03550_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08224_  (.A(\soc/cpu/_03550_ ),
    .B(\soc/cpu/_03538_ ),
    .Y(\soc/cpu/_03551_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_08225_  (.A(\soc/cpu/decoded_imm[7] ),
    .B(\soc/cpu/reg_pc[7] ),
    .X(\soc/cpu/_03552_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08226_  (.A(\soc/cpu/decoded_imm[7] ),
    .B(\soc/cpu/reg_pc[7] ),
    .Y(\soc/cpu/_03553_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08227_  (.A(\soc/cpu/_03552_ ),
    .B(\soc/cpu/_03553_ ),
    .Y(\soc/cpu/_03554_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08228_  (.A(\soc/cpu/_03551_ ),
    .B(\soc/cpu/_03554_ ),
    .Y(\soc/cpu/_03555_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08229_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03555_ ),
    .Y(\soc/cpu/_03556_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08230_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[39] ),
    .B1(\soc/cpu/count_instr[7] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[39] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03557_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08231_  (.A(\soc/cpu/count_cycle[7] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03558_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08232_  (.A(\soc/cpu/_03021_ ),
    .Y(\soc/cpu/_03559_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08233_  (.A1(\soc/cpu/irq_mask[7] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[7] ),
    .C1(\soc/cpu/_03559_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03560_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_08234_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03557_ ),
    .B1(\soc/cpu/_03558_ ),
    .C1(\soc/cpu/_03560_ ),
    .Y(\soc/cpu/_03561_ ));
 sky130_fd_sc_hd__nand2_4 \soc/cpu/_08235_  (.A(net413),
    .B(\soc/cpu/_03561_ ),
    .Y(\soc/cpu/_03562_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08236_  (.A1(\soc/cpu/pcpi_rs1 [1]),
    .A2(\soc/mem_rdata[15] ),
    .B1(\soc/cpu/_03461_ ),
    .Y(\soc/cpu/_03563_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08237_  (.A1(\soc/cpu/pcpi_rs1 [1]),
    .A2(\soc/cpu/_02360_ ),
    .B1(\soc/cpu/_03563_ ),
    .Y(\soc/cpu/_03564_ ));
 sky130_fd_sc_hd__a221o_2 \soc/cpu/_08238_  (.A1(\soc/mem_rdata[7] ),
    .A2(\soc/cpu/mem_la_wstrb [0]),
    .B1(\soc/cpu/_03428_ ),
    .B2(\soc/mem_rdata[23] ),
    .C1(\soc/cpu/_03564_ ),
    .X(\soc/cpu/_03565_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08239_  (.A1(\soc/cpu/irq_pending[7] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03565_ ),
    .B2(\soc/cpu/cpu_state[6] ),
    .C1(\soc/cpu/cpu_state[4] ),
    .C2(net835),
    .Y(\soc/cpu/_03566_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08240_  (.A1(\soc/cpu/_03556_ ),
    .A2(\soc/cpu/_03562_ ),
    .A3(\soc/cpu/_03566_ ),
    .B1(net131),
    .Y(\soc/cpu/_00188_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08241_  (.A(\soc/cpu/decoded_imm[8] ),
    .B(net840),
    .Y(\soc/cpu/_03567_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_08242_  (.A(\soc/cpu/decoded_imm[8] ),
    .B(\soc/cpu/reg_pc[8] ),
    .X(\soc/cpu/_03568_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08243_  (.A(\soc/cpu/_03567_ ),
    .B(\soc/cpu/_03568_ ),
    .Y(\soc/cpu/_03569_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/cpu/_08244_  (.A1(\soc/cpu/_03535_ ),
    .A2(\soc/cpu/_03536_ ),
    .B1(\soc/cpu/_03553_ ),
    .C1(\soc/cpu/_03550_ ),
    .Y(\soc/cpu/_03570_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08245_  (.A(\soc/cpu/_03552_ ),
    .B(\soc/cpu/_03570_ ),
    .X(\soc/cpu/_03571_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08246_  (.A(\soc/cpu/_03569_ ),
    .B(\soc/cpu/_03571_ ),
    .Y(\soc/cpu/_03572_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_08247_  (.A(\soc/cpu/_03569_ ),
    .B(\soc/cpu/_03571_ ),
    .X(\soc/cpu/_03573_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08248_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03572_ ),
    .C(\soc/cpu/_03573_ ),
    .Y(\soc/cpu/_03574_ ));
 sky130_fd_sc_hd__and2_4 \soc/cpu/_08249_  (.A(\soc/cpu/latched_is_lb ),
    .B(\soc/cpu/_03565_ ),
    .X(\soc/cpu/_03575_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_08251_  (.A(\soc/cpu/latched_is_lh ),
    .B(\soc/cpu/latched_is_lb ),
    .Y(\soc/cpu/_03577_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_08252_  (.A(\soc/cpu/latched_is_lh ),
    .B(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03578_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08253_  (.A1(\soc/cpu/mem_wordsize[2] ),
    .A2(\soc/mem_rdata[8] ),
    .B1(\soc/cpu/_02283_ ),
    .Y(\soc/cpu/_03579_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_08254_  (.A1(\soc/cpu/mem_wordsize[2] ),
    .A2(\soc/cpu/_03425_ ),
    .B1(\soc/cpu/_03578_ ),
    .C1(\soc/cpu/_03579_ ),
    .Y(\soc/cpu/_03580_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08255_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03580_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03581_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08256_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[8] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03582_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08257_  (.A1(\soc/cpu/irq_mask[8] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[8] ),
    .C1(net159),
    .Y(\soc/cpu/_03583_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08258_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[40] ),
    .B1(\soc/cpu/count_instr[8] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[40] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03584_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08259_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03584_ ),
    .Y(\soc/cpu/_03585_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08260_  (.A1(\soc/cpu/count_cycle[8] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03585_ ),
    .Y(\soc/cpu/_03586_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08261_  (.A1(\soc/cpu/_03582_ ),
    .A2(\soc/cpu/_03583_ ),
    .B1(\soc/cpu/_03586_ ),
    .Y(\soc/cpu/_03587_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08262_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [8]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[8] ),
    .C1(net414),
    .C2(\soc/cpu/_03587_ ),
    .Y(\soc/cpu/_03588_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08263_  (.A1(\soc/cpu/_03574_ ),
    .A2(\soc/cpu/_03581_ ),
    .A3(\soc/cpu/_03588_ ),
    .B1(net131),
    .Y(\soc/cpu/_00189_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08264_  (.A(net874),
    .B(\soc/cpu/reg_pc[9] ),
    .Y(\soc/cpu/_03589_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08265_  (.A(net874),
    .B(\soc/cpu/reg_pc[9] ),
    .Y(\soc/cpu/_03590_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08266_  (.A(\soc/cpu/_03590_ ),
    .Y(\soc/cpu/_03591_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08267_  (.A(\soc/cpu/_03589_ ),
    .B(\soc/cpu/_03591_ ),
    .Y(\soc/cpu/_03592_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08268_  (.A1(\soc/cpu/_03569_ ),
    .A2(\soc/cpu/_03571_ ),
    .B1(\soc/cpu/_03568_ ),
    .Y(\soc/cpu/_03593_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08269_  (.A(\soc/cpu/_03592_ ),
    .B(\soc/cpu/_03593_ ),
    .Y(\soc/cpu/_03594_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08270_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03594_ ),
    .Y(\soc/cpu/_03595_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_08271_  (.A(\soc/cpu/mem_wordsize[2] ),
    .SLEEP(\soc/cpu/_03439_ ),
    .X(\soc/cpu/_03596_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08272_  (.A1(\soc/mem_rdata[9] ),
    .A2(net157),
    .B1(\soc/cpu/_03596_ ),
    .Y(\soc/cpu/_03597_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08273_  (.A(\soc/cpu/_03578_ ),
    .B(\soc/cpu/_03597_ ),
    .Y(\soc/cpu/_03598_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08274_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03598_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03599_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08275_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[41] ),
    .B1(\soc/cpu/count_instr[9] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[41] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03600_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08276_  (.A(\soc/cpu/count_cycle[9] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03601_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08277_  (.A(\soc/cpu/_03045_ ),
    .Y(\soc/cpu/_03602_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08278_  (.A1(\soc/cpu/irq_mask[9] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[9] ),
    .C1(\soc/cpu/_03602_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03603_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08279_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03600_ ),
    .B1(\soc/cpu/_03601_ ),
    .C1(net119),
    .Y(\soc/cpu/_03604_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08280_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [9]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[9] ),
    .C1(net414),
    .C2(\soc/cpu/_03604_ ),
    .Y(\soc/cpu/_03605_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08281_  (.A1(\soc/cpu/_03595_ ),
    .A2(\soc/cpu/_03599_ ),
    .A3(\soc/cpu/_03605_ ),
    .B1(net131),
    .Y(\soc/cpu/_00190_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08282_  (.A(net872),
    .B(\soc/cpu/reg_pc[10] ),
    .Y(\soc/cpu/_03606_ ));
 sky130_fd_sc_hd__a311oi_2 \soc/cpu/_08283_  (.A1(\soc/cpu/_03552_ ),
    .A2(\soc/cpu/_03569_ ),
    .A3(\soc/cpu/_03570_ ),
    .B1(\soc/cpu/_03591_ ),
    .C1(\soc/cpu/_03568_ ),
    .Y(\soc/cpu/_03607_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08284_  (.A(\soc/cpu/_03589_ ),
    .B(\soc/cpu/_03607_ ),
    .Y(\soc/cpu/_03608_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08285_  (.A(\soc/cpu/_03606_ ),
    .B(\soc/cpu/_03608_ ),
    .Y(\soc/cpu/_03609_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08286_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03609_ ),
    .Y(\soc/cpu/_03610_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08287_  (.A1(\soc/mem_rdata[10] ),
    .A2(net157),
    .B1(\soc/cpu/_03460_ ),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_03611_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08288_  (.A(\soc/cpu/_03578_ ),
    .B(\soc/cpu/_03611_ ),
    .Y(\soc/cpu/_03612_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08289_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03612_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03613_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08291_  (.A1(\soc/cpu/irq_mask[10] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[10] ),
    .C1(net159),
    .X(\soc/cpu/_03615_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/cpu/_08292_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/cpuregs_rdata1[10] ),
    .A3(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_03615_ ),
    .Y(\soc/cpu/_03616_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08293_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[42] ),
    .B1(\soc/cpu/count_instr[10] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[42] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03617_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08294_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03617_ ),
    .Y(\soc/cpu/_03618_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08295_  (.A1(\soc/cpu/count_cycle[10] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03618_ ),
    .C1(net413),
    .Y(\soc/cpu/_03619_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08296_  (.A1(\soc/cpu/_03616_ ),
    .A2(\soc/cpu/_03619_ ),
    .B1(_074_),
    .Y(\soc/cpu/_03620_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_08297_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [10]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[10] ),
    .C1(\soc/cpu/_03620_ ),
    .Y(\soc/cpu/_03621_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08298_  (.A(\soc/cpu/_03610_ ),
    .B(\soc/cpu/_03613_ ),
    .C(\soc/cpu/_03621_ ),
    .Y(\soc/cpu/_00191_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08299_  (.A(\soc/cpu/decoded_imm[11] ),
    .B(\soc/cpu/reg_pc[11] ),
    .Y(\soc/cpu/_03622_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08300_  (.A(net872),
    .B(\soc/cpu/reg_pc[10] ),
    .Y(\soc/cpu/_03623_ ));
 sky130_fd_sc_hd__o31a_1 \soc/cpu/_08301_  (.A1(\soc/cpu/_03589_ ),
    .A2(\soc/cpu/_03606_ ),
    .A3(\soc/cpu/_03607_ ),
    .B1(\soc/cpu/_03623_ ),
    .X(\soc/cpu/_03624_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08302_  (.A(\soc/cpu/_03622_ ),
    .B(\soc/cpu/_03624_ ),
    .Y(\soc/cpu/_03625_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08303_  (.A(\soc/cpu/_03622_ ),
    .B(\soc/cpu/_03624_ ),
    .Y(\soc/cpu/_03626_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_08304_  (.A_N(\soc/cpu/_03625_ ),
    .B(\soc/cpu/_03626_ ),
    .C(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03627_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_08305_  (.A1(\soc/mem_rdata[11] ),
    .A2(net157),
    .B1(\soc/cpu/_03475_ ),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_03628_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08306_  (.A(\soc/cpu/_03578_ ),
    .B(\soc/cpu/_03628_ ),
    .Y(\soc/cpu/_03629_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08307_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03629_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03630_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08308_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[43] ),
    .B1(\soc/cpu/count_instr[11] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[43] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03631_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08309_  (.A(\soc/cpu/count_cycle[11] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03632_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08310_  (.A(\soc/cpu/_03068_ ),
    .Y(\soc/cpu/_03633_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08311_  (.A1(\soc/cpu/irq_mask[11] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[11] ),
    .C1(\soc/cpu/_03633_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03634_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08312_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03631_ ),
    .B1(\soc/cpu/_03632_ ),
    .C1(net118),
    .Y(\soc/cpu/_03635_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08313_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [11]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[11] ),
    .C1(net414),
    .C2(\soc/cpu/_03635_ ),
    .Y(\soc/cpu/_03636_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08314_  (.A1(\soc/cpu/_03627_ ),
    .A2(\soc/cpu/_03630_ ),
    .A3(\soc/cpu/_03636_ ),
    .B1(net131),
    .Y(\soc/cpu/_00192_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08315_  (.A(\soc/cpu/decoded_imm[11] ),
    .B(\soc/cpu/reg_pc[11] ),
    .X(\soc/cpu/_03637_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_08316_  (.A(net948),
    .B(\soc/cpu/reg_pc[12] ),
    .X(\soc/cpu/_03638_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08317_  (.A1(\soc/cpu/_03637_ ),
    .A2(\soc/cpu/_03625_ ),
    .B1(\soc/cpu/_03638_ ),
    .Y(\soc/cpu/_03639_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_08318_  (.A(\soc/cpu/_03637_ ),
    .B(\soc/cpu/_03625_ ),
    .C(\soc/cpu/_03638_ ),
    .X(\soc/cpu/_03640_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08319_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03639_ ),
    .C(\soc/cpu/_03640_ ),
    .Y(\soc/cpu/_03641_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_08320_  (.A1(\soc/mem_rdata[12] ),
    .A2(net157),
    .B1(\soc/cpu/_03504_ ),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_03642_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08321_  (.A(\soc/cpu/_03578_ ),
    .B(\soc/cpu/_03642_ ),
    .Y(\soc/cpu/_03643_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08322_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03643_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03644_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08323_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[44] ),
    .B1(\soc/cpu/count_instr[12] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[44] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03645_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08324_  (.A(\soc/cpu/count_cycle[12] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03646_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08325_  (.A(\soc/cpu/_03076_ ),
    .Y(\soc/cpu/_03647_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08326_  (.A1(\soc/cpu/irq_mask[12] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[12] ),
    .C1(\soc/cpu/_03647_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03648_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08327_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03645_ ),
    .B1(\soc/cpu/_03646_ ),
    .C1(net117),
    .Y(\soc/cpu/_03649_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08328_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [12]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[12] ),
    .C1(net414),
    .C2(\soc/cpu/_03649_ ),
    .Y(\soc/cpu/_03650_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08329_  (.A1(\soc/cpu/_03641_ ),
    .A2(\soc/cpu/_03644_ ),
    .A3(\soc/cpu/_03650_ ),
    .B1(net131),
    .Y(\soc/cpu/_00193_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08330_  (.A(\soc/cpu/decoded_imm[13] ),
    .B(\soc/cpu/reg_pc[13] ),
    .Y(\soc/cpu/_03651_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08331_  (.A(\soc/cpu/_03651_ ),
    .Y(\soc/cpu/_03652_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08332_  (.A(\soc/cpu/decoded_imm[13] ),
    .B(\soc/cpu/reg_pc[13] ),
    .Y(\soc/cpu/_03653_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08333_  (.A(\soc/cpu/_03652_ ),
    .B(\soc/cpu/_03653_ ),
    .Y(\soc/cpu/_03654_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08334_  (.A(\soc/cpu/decoded_imm[12] ),
    .B(\soc/cpu/reg_pc[12] ),
    .Y(\soc/cpu/_03655_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08335_  (.A(\soc/cpu/_03655_ ),
    .B(\soc/cpu/_03639_ ),
    .X(\soc/cpu/_03656_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08336_  (.A(\soc/cpu/_03654_ ),
    .B(\soc/cpu/_03656_ ),
    .Y(\soc/cpu/_03657_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_08337_  (.A1(\soc/cpu/_03654_ ),
    .A2(\soc/cpu/_03656_ ),
    .B1(\soc/cpu/_03657_ ),
    .C1(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03658_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_08338_  (.A1(\soc/mem_rdata[13] ),
    .A2(net157),
    .B1(\soc/cpu/_03514_ ),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_03659_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08339_  (.A(\soc/cpu/_03578_ ),
    .B(\soc/cpu/_03659_ ),
    .Y(\soc/cpu/_03660_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08340_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03660_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03661_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08341_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[45] ),
    .B1(\soc/cpu/count_instr[13] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[45] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03662_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08342_  (.A(\soc/cpu/count_cycle[13] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03663_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08343_  (.A(\soc/cpu/_03090_ ),
    .Y(\soc/cpu/_03664_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08344_  (.A1(\soc/cpu/irq_mask[13] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[13] ),
    .C1(\soc/cpu/_03664_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03665_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08345_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03662_ ),
    .B1(\soc/cpu/_03663_ ),
    .C1(net116),
    .Y(\soc/cpu/_03666_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08346_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [13]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[13] ),
    .C1(net414),
    .C2(\soc/cpu/_03666_ ),
    .Y(\soc/cpu/_03667_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08347_  (.A1(\soc/cpu/_03658_ ),
    .A2(\soc/cpu/_03661_ ),
    .A3(\soc/cpu/_03667_ ),
    .B1(net131),
    .Y(\soc/cpu/_00194_ ));
 sky130_fd_sc_hd__o2111ai_2 \soc/cpu/_08348_  (.A1(\soc/cpu/_03637_ ),
    .A2(\soc/cpu/_03625_ ),
    .B1(\soc/cpu/_03638_ ),
    .C1(\soc/cpu/_03652_ ),
    .D1(\soc/cpu/_03653_ ),
    .Y(\soc/cpu/_03668_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_08349_  (.A1(\soc/cpu/_03655_ ),
    .A2(\soc/cpu/_03651_ ),
    .B1(\soc/cpu/_03653_ ),
    .X(\soc/cpu/_03669_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08350_  (.A(\soc/cpu/decoded_imm[14] ),
    .B(\soc/cpu/reg_pc[14] ),
    .Y(\soc/cpu/_03670_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_08351_  (.A1(\soc/cpu/_03668_ ),
    .A2(\soc/cpu/_03669_ ),
    .B1(\soc/cpu/_03670_ ),
    .X(\soc/cpu/_03671_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08352_  (.A(\soc/cpu/_03668_ ),
    .B(\soc/cpu/_03670_ ),
    .C(\soc/cpu/_03669_ ),
    .Y(\soc/cpu/_03672_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08353_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03671_ ),
    .C(\soc/cpu/_03672_ ),
    .Y(\soc/cpu/_03673_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/_08354_  (.A1(\soc/mem_rdata[14] ),
    .A2(net157),
    .B1(\soc/cpu/_03546_ ),
    .B2(\soc/cpu/mem_wordsize[2] ),
    .Y(\soc/cpu/_03674_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08355_  (.A(\soc/cpu/_03578_ ),
    .B(\soc/cpu/_03674_ ),
    .Y(\soc/cpu/_03675_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08356_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03675_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03676_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08357_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[46] ),
    .B1(\soc/cpu/count_instr[14] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[46] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03677_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08358_  (.A1(\soc/cpu/count_cycle[14] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(net413),
    .Y(\soc/cpu/_03678_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08359_  (.A1(\soc/cpu/irq_mask[14] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[14] ),
    .C1(net159),
    .X(\soc/cpu/_03679_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/cpu/_08360_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/cpuregs_rdata1[14] ),
    .A3(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_03679_ ),
    .Y(\soc/cpu/_03680_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/cpu/_08361_  (.A1(\soc/cpu/_03414_ ),
    .A2(\soc/cpu/_03677_ ),
    .B1(\soc/cpu/_03678_ ),
    .C1(\soc/cpu/_03680_ ),
    .Y(\soc/cpu/_03681_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08362_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [14]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[14] ),
    .C1(\soc/cpu/_03681_ ),
    .Y(\soc/cpu/_03682_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08363_  (.A1(\soc/cpu/_03673_ ),
    .A2(\soc/cpu/_03676_ ),
    .A3(\soc/cpu/_03682_ ),
    .B1(net131),
    .Y(\soc/cpu/_00195_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08365_  (.A(\soc/cpu/decoded_imm[15] ),
    .B(\soc/cpu/reg_pc[15] ),
    .Y(\soc/cpu/_03684_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08366_  (.A(\soc/cpu/decoded_imm[15] ),
    .B(\soc/cpu/reg_pc[15] ),
    .Y(\soc/cpu/_03685_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_08367_  (.A(\soc/cpu/_03684_ ),
    .B_N(\soc/cpu/_03685_ ),
    .Y(\soc/cpu/_03686_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08368_  (.A(\soc/cpu/decoded_imm[14] ),
    .B(\soc/cpu/reg_pc[14] ),
    .Y(\soc/cpu/_03687_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08369_  (.A(\soc/cpu/_03687_ ),
    .B(\soc/cpu/_03671_ ),
    .X(\soc/cpu/_03688_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08370_  (.A(\soc/cpu/_03686_ ),
    .B(\soc/cpu/_03688_ ),
    .Y(\soc/cpu/_03689_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08371_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[15] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03690_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08372_  (.A1(\soc/cpu/irq_mask[15] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[15] ),
    .C1(net159),
    .Y(\soc/cpu/_03691_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08373_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[47] ),
    .B1(\soc/cpu/count_instr[15] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[47] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03692_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08374_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03692_ ),
    .Y(\soc/cpu/_03693_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08375_  (.A1(\soc/cpu/count_cycle[15] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03693_ ),
    .Y(\soc/cpu/_03694_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08376_  (.A1(\soc/cpu/_03690_ ),
    .A2(\soc/cpu/_03691_ ),
    .B1(\soc/cpu/_03694_ ),
    .Y(\soc/cpu/_03695_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08377_  (.A(\soc/mem_rdata[15] ),
    .B(\soc/cpu/_02282_ ),
    .C(\soc/cpu/_02283_ ),
    .Y(\soc/cpu/_03696_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_08378_  (.A1(\soc/cpu/_02360_ ),
    .A2(\soc/cpu/_02282_ ),
    .B1(\soc/cpu/_03696_ ),
    .X(\soc/cpu/_03697_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_08379_  (.A(\soc/cpu/latched_is_lh ),
    .SLEEP(\soc/cpu/_03697_ ),
    .X(\soc/cpu/_03698_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_08380_  (.A1(\soc/cpu/_03575_ ),
    .A2(\soc/cpu/_03577_ ),
    .A3(\soc/cpu/_03698_ ),
    .B1(\soc/cpu/cpu_state[6] ),
    .Y(\soc/cpu/_03699_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08381_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03697_ ),
    .B1(\soc/cpu/_03699_ ),
    .Y(\soc/cpu/_03700_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08382_  (.A1(\soc/cpu/irq_pending[15] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03695_ ),
    .B2(net414),
    .C1(\soc/cpu/_03700_ ),
    .X(\soc/cpu/_03701_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08383_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [15]),
    .B1(\soc/cpu/_03689_ ),
    .B2(\soc/cpu/cpu_state[3] ),
    .C1(\soc/cpu/_03701_ ),
    .Y(\soc/cpu/_03702_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08384_  (.A(net131),
    .B(\soc/cpu/_03702_ ),
    .Y(\soc/cpu/_00196_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08385_  (.A(\soc/cpu/decoded_imm[16] ),
    .B(\soc/cpu/reg_pc[16] ),
    .Y(\soc/cpu/_03703_ ));
 sky130_fd_sc_hd__a311o_2 \soc/cpu/_08386_  (.A1(\soc/cpu/_03687_ ),
    .A2(\soc/cpu/_03671_ ),
    .A3(\soc/cpu/_03685_ ),
    .B1(\soc/cpu/_03703_ ),
    .C1(\soc/cpu/_03684_ ),
    .X(\soc/cpu/_03704_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_08387_  (.A1(\soc/cpu/_03684_ ),
    .A2(\soc/cpu/_03688_ ),
    .B1(\soc/cpu/_03703_ ),
    .C1(\soc/cpu/_03685_ ),
    .Y(\soc/cpu/_03705_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08390_  (.A1(\soc/mem_rdata[16] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03708_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08391_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[16] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03709_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08392_  (.A1(\soc/cpu/irq_mask[16] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[16] ),
    .C1(net159),
    .Y(\soc/cpu/_03710_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08393_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[48] ),
    .B1(\soc/cpu/count_instr[16] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[48] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03711_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08394_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03711_ ),
    .Y(\soc/cpu/_03712_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08395_  (.A1(\soc/cpu/count_cycle[16] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03712_ ),
    .Y(\soc/cpu/_03713_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08396_  (.A1(\soc/cpu/_03709_ ),
    .A2(\soc/cpu/_03710_ ),
    .B1(\soc/cpu/_03713_ ),
    .Y(\soc/cpu/_03714_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08397_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [16]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[16] ),
    .C1(net414),
    .C2(\soc/cpu/_03714_ ),
    .Y(\soc/cpu/_03715_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08398_  (.A1(net53),
    .A2(\soc/cpu/_03708_ ),
    .B1(\soc/cpu/_03715_ ),
    .Y(\soc/cpu/_03716_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08399_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03704_ ),
    .A3(\soc/cpu/_03705_ ),
    .B1(\soc/cpu/_03716_ ),
    .Y(\soc/cpu/_03717_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08400_  (.A(net131),
    .B(\soc/cpu/_03717_ ),
    .Y(\soc/cpu/_00197_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_08401_  (.A(\soc/cpu/decoded_imm[17] ),
    .B(\soc/cpu/reg_pc[17] ),
    .Y(\soc/cpu/_03718_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08402_  (.A(\soc/cpu/decoded_imm[17] ),
    .B(\soc/cpu/reg_pc[17] ),
    .X(\soc/cpu/_03719_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08403_  (.A(\soc/cpu/decoded_imm[16] ),
    .B(\soc/cpu/reg_pc[16] ),
    .Y(\soc/cpu/_03720_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08404_  (.A(\soc/cpu/_03720_ ),
    .B(\soc/cpu/_03704_ ),
    .X(\soc/cpu/_03721_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08405_  (.A1(\soc/cpu/_03718_ ),
    .A2(\soc/cpu/_03719_ ),
    .B1(\soc/cpu/_03721_ ),
    .Y(\soc/cpu/_03722_ ));
 sky130_fd_sc_hd__o311ai_1 \soc/cpu/_08406_  (.A1(\soc/cpu/_03718_ ),
    .A2(\soc/cpu/_03719_ ),
    .A3(\soc/cpu/_03721_ ),
    .B1(\soc/cpu/_03722_ ),
    .C1(\soc/cpu/cpu_state[3] ),
    .Y(\soc/cpu/_03723_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08407_  (.A(\soc/cpu/cpu_state[4] ),
    .B(net888),
    .Y(\soc/cpu/_03724_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08408_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[17] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03725_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08409_  (.A1(\soc/cpu/irq_mask[17] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[17] ),
    .C1(net159),
    .Y(\soc/cpu/_03726_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08410_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[49] ),
    .B1(\soc/cpu/count_instr[17] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[49] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03727_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08411_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03727_ ),
    .Y(\soc/cpu/_03728_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08412_  (.A1(\soc/cpu/count_cycle[17] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03728_ ),
    .Y(\soc/cpu/_03729_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08413_  (.A1(\soc/cpu/_03725_ ),
    .A2(\soc/cpu/_03726_ ),
    .B1(\soc/cpu/_03729_ ),
    .Y(\soc/cpu/_03730_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08414_  (.A(\soc/mem_rdata[17] ),
    .B(net157),
    .Y(\soc/cpu/_03731_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08415_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03731_ ),
    .B1(\soc/cpu/_03699_ ),
    .Y(\soc/cpu/_03732_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_08416_  (.A1(\soc/cpu/irq_pending[17] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03730_ ),
    .B2(net414),
    .C1(\soc/cpu/_03732_ ),
    .Y(\soc/cpu/_03733_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08417_  (.A1(\soc/cpu/_03723_ ),
    .A2(\soc/cpu/_03724_ ),
    .A3(\soc/cpu/_03733_ ),
    .B1(net131),
    .Y(\soc/cpu/_00198_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_08418_  (.A(\soc/cpu/decoded_imm[18] ),
    .B(\soc/cpu/reg_pc[18] ),
    .Y(\soc/cpu/_03734_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08419_  (.A(\soc/cpu/decoded_imm[17] ),
    .B(\soc/cpu/reg_pc[17] ),
    .Y(\soc/cpu/_03735_ ));
 sky130_fd_sc_hd__o211a_1 \soc/cpu/_08420_  (.A1(\soc/cpu/_03718_ ),
    .A2(\soc/cpu/_03721_ ),
    .B1(\soc/cpu/_03734_ ),
    .C1(\soc/cpu/_03735_ ),
    .X(\soc/cpu/_03736_ ));
 sky130_fd_sc_hd__a311oi_4 \soc/cpu/_08421_  (.A1(\soc/cpu/_03720_ ),
    .A2(\soc/cpu/_03704_ ),
    .A3(\soc/cpu/_03735_ ),
    .B1(\soc/cpu/_03734_ ),
    .C1(\soc/cpu/_03718_ ),
    .Y(\soc/cpu/_03737_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08422_  (.A(\soc/mem_rdata[18] ),
    .B(net157),
    .Y(\soc/cpu/_03738_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08423_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03738_ ),
    .B1(\soc/cpu/_03699_ ),
    .Y(\soc/cpu/_03739_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08424_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[50] ),
    .B1(\soc/cpu/count_instr[18] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[50] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03740_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08425_  (.A1(\soc/cpu/count_cycle[18] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(net413),
    .Y(\soc/cpu/_03741_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08426_  (.A1(\soc/cpu/irq_mask[18] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[18] ),
    .C1(\soc/cpu/_00872_ ),
    .X(\soc/cpu/_03742_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/cpu/_08427_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/cpuregs_rdata1[18] ),
    .A3(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_03742_ ),
    .Y(\soc/cpu/_03743_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/cpu/_08428_  (.A1(\soc/cpu/_03414_ ),
    .A2(\soc/cpu/_03740_ ),
    .B1(\soc/cpu/_03741_ ),
    .C1(\soc/cpu/_03743_ ),
    .Y(\soc/cpu/_03744_ ));
 sky130_fd_sc_hd__a221o_2 \soc/cpu/_08429_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [18]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[18] ),
    .C1(\soc/cpu/_03744_ ),
    .X(\soc/cpu/_03745_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08430_  (.A(\soc/cpu/_03739_ ),
    .B(\soc/cpu/_03745_ ),
    .Y(\soc/cpu/_03746_ ));
 sky130_fd_sc_hd__o31a_1 \soc/cpu/_08431_  (.A1(\soc/cpu/_00940_ ),
    .A2(\soc/cpu/_03736_ ),
    .A3(\soc/cpu/_03737_ ),
    .B1(\soc/cpu/_03746_ ),
    .X(\soc/cpu/_03747_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08432_  (.A(net131),
    .B(\soc/cpu/_03747_ ),
    .Y(\soc/cpu/_00199_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08433_  (.A(\soc/cpu/decoded_imm[18] ),
    .B(\soc/cpu/reg_pc[18] ),
    .Y(\soc/cpu/_03748_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08434_  (.A(\soc/cpu/_03748_ ),
    .Y(\soc/cpu/_03749_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08435_  (.A(\soc/cpu/decoded_imm[19] ),
    .B(\soc/cpu/reg_pc[19] ),
    .Y(\soc/cpu/_03750_ ));
 sky130_fd_sc_hd__o21bai_2 \soc/cpu/_08436_  (.A1(\soc/cpu/_03749_ ),
    .A2(\soc/cpu/_03737_ ),
    .B1_N(\soc/cpu/_03750_ ),
    .Y(\soc/cpu/_03751_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08437_  (.A(\soc/cpu/_03749_ ),
    .B(\soc/cpu/_03737_ ),
    .Y(\soc/cpu/_03752_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08438_  (.A1(\soc/cpu/_03750_ ),
    .A2(\soc/cpu/_03752_ ),
    .B1(\soc/cpu/_00940_ ),
    .Y(\soc/cpu/_03753_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08439_  (.A(\soc/cpu/_03751_ ),
    .B(\soc/cpu/_03753_ ),
    .Y(\soc/cpu/_03754_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08440_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/pcpi_rs1 [19]),
    .Y(\soc/cpu/_03755_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08441_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[19] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03756_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08442_  (.A1(\soc/cpu/irq_mask[19] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[19] ),
    .C1(net159),
    .Y(\soc/cpu/_03757_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08443_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[51] ),
    .B1(\soc/cpu/count_instr[19] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[51] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03758_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08444_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03758_ ),
    .Y(\soc/cpu/_03759_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08445_  (.A1(\soc/cpu/count_cycle[19] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03759_ ),
    .Y(\soc/cpu/_03760_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08446_  (.A1(\soc/cpu/_03756_ ),
    .A2(\soc/cpu/_03757_ ),
    .B1(\soc/cpu/_03760_ ),
    .Y(\soc/cpu/_03761_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08447_  (.A(\soc/mem_rdata[19] ),
    .B(net157),
    .Y(\soc/cpu/_03762_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08448_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03762_ ),
    .B1(net54),
    .Y(\soc/cpu/_03763_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_08449_  (.A1(\soc/cpu/irq_pending[19] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03761_ ),
    .B2(net414),
    .C1(\soc/cpu/_03763_ ),
    .Y(\soc/cpu/_03764_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08450_  (.A1(\soc/cpu/_03754_ ),
    .A2(\soc/cpu/_03755_ ),
    .A3(\soc/cpu/_03764_ ),
    .B1(net131),
    .Y(\soc/cpu/_00200_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08451_  (.A(\soc/cpu/decoded_imm[19] ),
    .B(\soc/cpu/reg_pc[19] ),
    .Y(\soc/cpu/_03765_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08452_  (.A(\soc/cpu/decoded_imm[20] ),
    .B(\soc/cpu/reg_pc[20] ),
    .Y(\soc/cpu/_03766_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08453_  (.A(\soc/cpu/decoded_imm[20] ),
    .B(\soc/cpu/reg_pc[20] ),
    .X(\soc/cpu/_03767_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/_08454_  (.A1(\soc/cpu/_03765_ ),
    .A2(\soc/cpu/_03751_ ),
    .B1(\soc/cpu/_03766_ ),
    .C1(\soc/cpu/_03767_ ),
    .X(\soc/cpu/_03768_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_08455_  (.A1(\soc/cpu/_03766_ ),
    .A2(\soc/cpu/_03767_ ),
    .B1(\soc/cpu/_03765_ ),
    .C1(\soc/cpu/_03751_ ),
    .Y(\soc/cpu/_03769_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08456_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03768_ ),
    .C(\soc/cpu/_03769_ ),
    .Y(\soc/cpu/_03770_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08457_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/pcpi_rs1 [20]),
    .Y(\soc/cpu/_03771_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08458_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[20] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03772_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08459_  (.A1(\soc/cpu/irq_mask[20] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[20] ),
    .C1(net159),
    .Y(\soc/cpu/_03773_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08460_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[52] ),
    .B1(\soc/cpu/count_instr[20] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[52] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03774_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08461_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03774_ ),
    .Y(\soc/cpu/_03775_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08462_  (.A1(\soc/cpu/count_cycle[20] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03775_ ),
    .Y(\soc/cpu/_03776_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08463_  (.A1(\soc/cpu/_03772_ ),
    .A2(\soc/cpu/_03773_ ),
    .B1(\soc/cpu/_03776_ ),
    .Y(\soc/cpu/_03777_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08464_  (.A(\soc/mem_rdata[20] ),
    .B(net157),
    .Y(\soc/cpu/_03778_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08465_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03778_ ),
    .B1(\soc/cpu/_03699_ ),
    .Y(\soc/cpu/_03779_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_08466_  (.A1(\soc/cpu/irq_pending[20] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03777_ ),
    .B2(net414),
    .C1(\soc/cpu/_03779_ ),
    .Y(\soc/cpu/_03780_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08467_  (.A1(\soc/cpu/_03770_ ),
    .A2(\soc/cpu/_03771_ ),
    .A3(\soc/cpu/_03780_ ),
    .B1(net131),
    .Y(\soc/cpu/_00201_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08468_  (.A(\soc/cpu/decoded_imm[20] ),
    .B(\soc/cpu/reg_pc[20] ),
    .Y(\soc/cpu/_03781_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08469_  (.A(\soc/cpu/decoded_imm[21] ),
    .B(\soc/cpu/reg_pc[21] ),
    .Y(\soc/cpu/_03782_ ));
 sky130_fd_sc_hd__a2111o_1 \soc/cpu/_08470_  (.A1(\soc/cpu/_03765_ ),
    .A2(\soc/cpu/_03751_ ),
    .B1(\soc/cpu/_03766_ ),
    .C1(\soc/cpu/_03767_ ),
    .D1(\soc/cpu/_03782_ ),
    .X(\soc/cpu/_03783_ ));
 sky130_fd_sc_hd__or2_1 \soc/cpu/_08471_  (.A(\soc/cpu/_03781_ ),
    .B(\soc/cpu/_03782_ ),
    .X(\soc/cpu/_03784_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08472_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03783_ ),
    .C(\soc/cpu/_03784_ ),
    .Y(\soc/cpu/_03785_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_08473_  (.A1(\soc/cpu/_03781_ ),
    .A2(\soc/cpu/_03768_ ),
    .A3(\soc/cpu/_03782_ ),
    .B1(\soc/cpu/_03785_ ),
    .Y(\soc/cpu/_03786_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08474_  (.A(\soc/mem_rdata[21] ),
    .B(net157),
    .Y(\soc/cpu/_03787_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08475_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03787_ ),
    .B1(net54),
    .Y(\soc/cpu/_03788_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08476_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[53] ),
    .B1(\soc/cpu/count_instr[21] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[53] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03789_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08477_  (.A1(\soc/cpu/count_cycle[21] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(net413),
    .Y(\soc/cpu/_03790_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08478_  (.A1(\soc/cpu/irq_mask[21] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[21] ),
    .C1(\soc/cpu/_00872_ ),
    .X(\soc/cpu/_03791_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/cpu/_08479_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/cpuregs_rdata1[21] ),
    .A3(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_03791_ ),
    .Y(\soc/cpu/_03792_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/cpu/_08480_  (.A1(\soc/cpu/_03414_ ),
    .A2(\soc/cpu/_03789_ ),
    .B1(\soc/cpu/_03790_ ),
    .C1(\soc/cpu/_03792_ ),
    .Y(\soc/cpu/_03793_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08481_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [21]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[21] ),
    .C1(\soc/cpu/_03793_ ),
    .X(\soc/cpu/_03794_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08482_  (.A(\soc/cpu/_03786_ ),
    .B(\soc/cpu/_03788_ ),
    .C(\soc/cpu/_03794_ ),
    .Y(\soc/cpu/_03795_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08483_  (.A(net131),
    .B(\soc/cpu/_03795_ ),
    .Y(\soc/cpu/_00202_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08484_  (.A(\soc/cpu/decoded_imm[22] ),
    .B(\soc/cpu/reg_pc[22] ),
    .Y(\soc/cpu/_03796_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08485_  (.A(\soc/cpu/decoded_imm[21] ),
    .B(\soc/cpu/reg_pc[21] ),
    .Y(\soc/cpu/_03797_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08486_  (.A(\soc/cpu/_03797_ ),
    .B(\soc/cpu/_03783_ ),
    .C(\soc/cpu/_03784_ ),
    .Y(\soc/cpu/_03798_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08487_  (.A(\soc/cpu/_03796_ ),
    .B(\soc/cpu/_03798_ ),
    .Y(\soc/cpu/_03799_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08488_  (.A1(\soc/mem_rdata[22] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03800_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08489_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[22] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03801_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08490_  (.A1(\soc/cpu/irq_mask[22] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[22] ),
    .C1(net159),
    .Y(\soc/cpu/_03802_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08491_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[54] ),
    .B1(\soc/cpu/count_instr[22] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[54] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03803_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08492_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03803_ ),
    .Y(\soc/cpu/_03804_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08493_  (.A1(\soc/cpu/count_cycle[22] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03804_ ),
    .Y(\soc/cpu/_03805_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08494_  (.A1(\soc/cpu/_03801_ ),
    .A2(\soc/cpu/_03802_ ),
    .B1(\soc/cpu/_03805_ ),
    .Y(\soc/cpu/_03806_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08495_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [22]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[22] ),
    .C1(net414),
    .C2(\soc/cpu/_03806_ ),
    .Y(\soc/cpu/_03807_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08496_  (.A1(net53),
    .A2(\soc/cpu/_03800_ ),
    .B1(\soc/cpu/_03807_ ),
    .Y(\soc/cpu/_03808_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08497_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03799_ ),
    .B1(\soc/cpu/_03808_ ),
    .Y(\soc/cpu/_03809_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08498_  (.A(net131),
    .B(\soc/cpu/_03809_ ),
    .Y(\soc/cpu/_00203_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08499_  (.A(\soc/cpu/decoded_imm[23] ),
    .B(\soc/cpu/reg_pc[23] ),
    .Y(\soc/cpu/_03810_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08500_  (.A1(\soc/cpu/_03797_ ),
    .A2(\soc/cpu/_03783_ ),
    .A3(\soc/cpu/_03784_ ),
    .B1(\soc/cpu/_03796_ ),
    .Y(\soc/cpu/_03811_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08501_  (.A1(\soc/cpu/decoded_imm[22] ),
    .A2(\soc/cpu/reg_pc[22] ),
    .B1(\soc/cpu/_03811_ ),
    .Y(\soc/cpu/_03812_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08502_  (.A(\soc/cpu/decoded_imm[22] ),
    .B(\soc/cpu/reg_pc[22] ),
    .Y(\soc/cpu/_03813_ ));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_08503_  (.A(\soc/cpu/_03813_ ),
    .B(\soc/cpu/_03810_ ),
    .X(\soc/cpu/_03814_ ));
 sky130_fd_sc_hd__a311o_2 \soc/cpu/_08504_  (.A1(\soc/cpu/_03797_ ),
    .A2(\soc/cpu/_03783_ ),
    .A3(\soc/cpu/_03784_ ),
    .B1(\soc/cpu/_03796_ ),
    .C1(\soc/cpu/_03810_ ),
    .X(\soc/cpu/_03815_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08505_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03814_ ),
    .C(\soc/cpu/_03815_ ),
    .Y(\soc/cpu/_03816_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08506_  (.A1(\soc/cpu/_03810_ ),
    .A2(\soc/cpu/_03812_ ),
    .B1(\soc/cpu/_03816_ ),
    .Y(\soc/cpu/_03817_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08507_  (.A1(\soc/mem_rdata[23] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03818_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08508_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[23] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03819_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08509_  (.A1(\soc/cpu/irq_mask[23] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[23] ),
    .C1(net159),
    .Y(\soc/cpu/_03820_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08510_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[55] ),
    .B1(\soc/cpu/count_instr[23] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[55] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03821_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08511_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03821_ ),
    .Y(\soc/cpu/_03822_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08512_  (.A1(\soc/cpu/count_cycle[23] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03822_ ),
    .Y(\soc/cpu/_03823_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08513_  (.A1(\soc/cpu/_03819_ ),
    .A2(\soc/cpu/_03820_ ),
    .B1(\soc/cpu/_03823_ ),
    .Y(\soc/cpu/_03824_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08514_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [23]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[23] ),
    .C1(net414),
    .C2(\soc/cpu/_03824_ ),
    .Y(\soc/cpu/_03825_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08515_  (.A1(net53),
    .A2(\soc/cpu/_03818_ ),
    .B1(\soc/cpu/_03825_ ),
    .Y(\soc/cpu/_03826_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_08516_  (.A1(\soc/cpu/_03817_ ),
    .A2(\soc/cpu/_03826_ ),
    .B1(_074_),
    .X(\soc/cpu/_00204_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08517_  (.A(\soc/cpu/decoded_imm[23] ),
    .B(\soc/cpu/reg_pc[23] ),
    .Y(\soc/cpu/_03827_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_08518_  (.A(\soc/cpu/decoded_imm[24] ),
    .B(\soc/cpu/reg_pc[24] ),
    .Y(\soc/cpu/_03828_ ));
 sky130_fd_sc_hd__a31o_1 \soc/cpu/_08519_  (.A1(\soc/cpu/_03827_ ),
    .A2(\soc/cpu/_03814_ ),
    .A3(\soc/cpu/_03815_ ),
    .B1(\soc/cpu/_03828_ ),
    .X(\soc/cpu/_03829_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08520_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03829_ ),
    .Y(\soc/cpu/_03830_ ));
 sky130_fd_sc_hd__a41oi_4 \soc/cpu/_08521_  (.A1(\soc/cpu/_03827_ ),
    .A2(\soc/cpu/_03814_ ),
    .A3(\soc/cpu/_03815_ ),
    .A4(\soc/cpu/_03828_ ),
    .B1(\soc/cpu/_03830_ ),
    .Y(\soc/cpu/_03831_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08522_  (.A(\soc/mem_rdata[24] ),
    .B(net157),
    .Y(\soc/cpu/_03832_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08523_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03832_ ),
    .B1(net54),
    .Y(\soc/cpu/_03833_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08524_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[56] ),
    .B1(\soc/cpu/count_instr[24] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[56] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03834_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08525_  (.A1(\soc/cpu/count_cycle[24] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(net413),
    .Y(\soc/cpu/_03835_ ));
 sky130_fd_sc_hd__a221o_2 \soc/cpu/_08526_  (.A1(\soc/cpu/irq_mask[24] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[24] ),
    .C1(net159),
    .X(\soc/cpu/_03836_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_08527_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/cpuregs_rdata1[24] ),
    .A3(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_03836_ ),
    .Y(\soc/cpu/_03837_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/cpu/_08528_  (.A1(\soc/cpu/_03414_ ),
    .A2(\soc/cpu/_03834_ ),
    .B1(\soc/cpu/_03835_ ),
    .C1(\soc/cpu/_03837_ ),
    .Y(\soc/cpu/_03838_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08529_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [24]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[24] ),
    .C1(\soc/cpu/_03838_ ),
    .X(\soc/cpu/_03839_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08530_  (.A(\soc/cpu/_03831_ ),
    .B(\soc/cpu/_03833_ ),
    .C(\soc/cpu/_03839_ ),
    .Y(\soc/cpu/_03840_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08531_  (.A(net131),
    .B(\soc/cpu/_03840_ ),
    .Y(\soc/cpu/_00205_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08532_  (.A(\soc/cpu/decoded_imm[24] ),
    .B(\soc/cpu/reg_pc[24] ),
    .Y(\soc/cpu/_03841_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08533_  (.A(\soc/cpu/_03841_ ),
    .B(\soc/cpu/_03829_ ),
    .X(\soc/cpu/_03842_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08534_  (.A(\soc/cpu/decoded_imm[25] ),
    .B(\soc/cpu/reg_pc[25] ),
    .Y(\soc/cpu/_03843_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08535_  (.A(\soc/cpu/decoded_imm[25] ),
    .B(\soc/cpu/reg_pc[25] ),
    .Y(\soc/cpu/_03844_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_08536_  (.A(\soc/cpu/_03843_ ),
    .B_N(\soc/cpu/_03844_ ),
    .Y(\soc/cpu/_03845_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08537_  (.A(\soc/cpu/_03842_ ),
    .B(\soc/cpu/_03845_ ),
    .Y(\soc/cpu/_03846_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08538_  (.A1(\soc/mem_rdata[25] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03847_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08539_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[57] ),
    .B1(\soc/cpu/count_instr[25] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[57] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03848_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08540_  (.A(\soc/cpu/count_cycle[25] ),
    .B(\soc/cpu/_00874_ ),
    .Y(\soc/cpu/_03849_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_08541_  (.A(\soc/cpu/_03223_ ),
    .Y(\soc/cpu/_03850_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08542_  (.A1(\soc/cpu/irq_mask[25] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[25] ),
    .C1(\soc/cpu/_03850_ ),
    .C2(\soc/cpu/instr_retirq ),
    .Y(\soc/cpu/_03851_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/cpu/_08543_  (.A1(\soc/cpu/_03446_ ),
    .A2(\soc/cpu/_03848_ ),
    .B1(\soc/cpu/_03849_ ),
    .C1(net115),
    .Y(\soc/cpu/_03852_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08544_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [25]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[25] ),
    .C1(net414),
    .C2(\soc/cpu/_03852_ ),
    .Y(\soc/cpu/_03853_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08545_  (.A1(net53),
    .A2(\soc/cpu/_03847_ ),
    .B1(\soc/cpu/_03853_ ),
    .Y(\soc/cpu/_03854_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08546_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03846_ ),
    .B1(\soc/cpu/_03854_ ),
    .Y(\soc/cpu/_03855_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08547_  (.A(net131),
    .B(\soc/cpu/_03855_ ),
    .Y(\soc/cpu/_00206_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08548_  (.A(\soc/cpu/decoded_imm[26] ),
    .B(\soc/cpu/reg_pc[26] ),
    .Y(\soc/cpu/_03856_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08549_  (.A1(\soc/cpu/_03842_ ),
    .A2(\soc/cpu/_03844_ ),
    .B1(\soc/cpu/_03843_ ),
    .Y(\soc/cpu/_03857_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08550_  (.A(\soc/cpu/_03856_ ),
    .B(\soc/cpu/_03857_ ),
    .Y(\soc/cpu/_03858_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08551_  (.A1(\soc/mem_rdata[26] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03859_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08552_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[26] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03860_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08553_  (.A1(\soc/cpu/irq_mask[26] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[26] ),
    .C1(net159),
    .Y(\soc/cpu/_03861_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08554_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[58] ),
    .B1(\soc/cpu/count_instr[26] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[58] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03862_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08555_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03862_ ),
    .Y(\soc/cpu/_03863_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08556_  (.A1(\soc/cpu/count_cycle[26] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03863_ ),
    .Y(\soc/cpu/_03864_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08557_  (.A1(\soc/cpu/_03860_ ),
    .A2(\soc/cpu/_03861_ ),
    .B1(\soc/cpu/_03864_ ),
    .Y(\soc/cpu/_03865_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08558_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [26]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[26] ),
    .C1(net414),
    .C2(\soc/cpu/_03865_ ),
    .Y(\soc/cpu/_03866_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08559_  (.A1(net53),
    .A2(\soc/cpu/_03859_ ),
    .B1(\soc/cpu/_03866_ ),
    .Y(\soc/cpu/_03867_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08560_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03858_ ),
    .B1(\soc/cpu/_03867_ ),
    .Y(\soc/cpu/_03868_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08561_  (.A(net131),
    .B(\soc/cpu/_03868_ ),
    .Y(\soc/cpu/_00207_ ));
 sky130_fd_sc_hd__a311oi_2 \soc/cpu/_08562_  (.A1(\soc/cpu/_03841_ ),
    .A2(\soc/cpu/_03829_ ),
    .A3(\soc/cpu/_03844_ ),
    .B1(\soc/cpu/_03856_ ),
    .C1(\soc/cpu/_03843_ ),
    .Y(\soc/cpu/_03869_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08563_  (.A1(\soc/cpu/decoded_imm[26] ),
    .A2(\soc/cpu/reg_pc[26] ),
    .B1(\soc/cpu/_03869_ ),
    .Y(\soc/cpu/_03870_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08564_  (.A(\soc/cpu/decoded_imm[27] ),
    .B(\soc/cpu/reg_pc[27] ),
    .Y(\soc/cpu/_03871_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08565_  (.A(\soc/cpu/decoded_imm[27] ),
    .B(\soc/cpu/reg_pc[27] ),
    .Y(\soc/cpu/_03872_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_08566_  (.A(\soc/cpu/_03871_ ),
    .B_N(\soc/cpu/_03872_ ),
    .Y(\soc/cpu/_03873_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08567_  (.A(\soc/cpu/_03870_ ),
    .B(\soc/cpu/_03873_ ),
    .Y(\soc/cpu/_03874_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08568_  (.A1(\soc/mem_rdata[27] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03875_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08569_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[27] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03876_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08570_  (.A1(\soc/cpu/irq_mask[27] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[27] ),
    .C1(net159),
    .Y(\soc/cpu/_03877_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08571_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[59] ),
    .B1(\soc/cpu/count_instr[27] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[59] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03878_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08572_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03878_ ),
    .Y(\soc/cpu/_03879_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08573_  (.A1(\soc/cpu/count_cycle[27] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03879_ ),
    .Y(\soc/cpu/_03880_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08574_  (.A1(\soc/cpu/_03876_ ),
    .A2(\soc/cpu/_03877_ ),
    .B1(\soc/cpu/_03880_ ),
    .Y(\soc/cpu/_03881_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08575_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [27]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[27] ),
    .C1(net414),
    .C2(\soc/cpu/_03881_ ),
    .Y(\soc/cpu/_03882_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08576_  (.A1(net53),
    .A2(\soc/cpu/_03875_ ),
    .B1(\soc/cpu/_03882_ ),
    .Y(\soc/cpu/_03883_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08577_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03874_ ),
    .B1(\soc/cpu/_03883_ ),
    .Y(\soc/cpu/_03884_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08578_  (.A(net131),
    .B(\soc/cpu/_03884_ ),
    .Y(\soc/cpu/_00208_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08579_  (.A(\soc/cpu/decoded_imm[28] ),
    .B(\soc/cpu/reg_pc[28] ),
    .Y(\soc/cpu/_03885_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08580_  (.A(\soc/cpu/decoded_imm[28] ),
    .B(\soc/cpu/reg_pc[28] ),
    .X(\soc/cpu/_03886_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08581_  (.A(\soc/cpu/_03885_ ),
    .B(\soc/cpu/_03886_ ),
    .Y(\soc/cpu/_03887_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08582_  (.A1(\soc/cpu/_03870_ ),
    .A2(\soc/cpu/_03872_ ),
    .B1(\soc/cpu/_03871_ ),
    .Y(\soc/cpu/_03888_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_08583_  (.A(\soc/cpu/_03887_ ),
    .B(\soc/cpu/_03888_ ),
    .X(\soc/cpu/_03889_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08584_  (.A1(\soc/mem_rdata[28] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03890_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08585_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[28] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03891_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08586_  (.A1(\soc/cpu/irq_mask[28] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[28] ),
    .C1(\soc/cpu/_00872_ ),
    .Y(\soc/cpu/_03892_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08587_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[60] ),
    .B1(\soc/cpu/count_instr[28] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[60] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03893_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08588_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03893_ ),
    .Y(\soc/cpu/_03894_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08589_  (.A1(\soc/cpu/count_cycle[28] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03894_ ),
    .Y(\soc/cpu/_03895_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08590_  (.A1(\soc/cpu/_03891_ ),
    .A2(\soc/cpu/_03892_ ),
    .B1(\soc/cpu/_03895_ ),
    .Y(\soc/cpu/_03896_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08591_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [28]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[28] ),
    .C1(net414),
    .C2(\soc/cpu/_03896_ ),
    .Y(\soc/cpu/_03897_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08592_  (.A1(net53),
    .A2(\soc/cpu/_03890_ ),
    .B1(\soc/cpu/_03897_ ),
    .Y(\soc/cpu/_03898_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08593_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03889_ ),
    .B1(\soc/cpu/_03898_ ),
    .Y(\soc/cpu/_03899_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08594_  (.A(net131),
    .B(\soc/cpu/_03899_ ),
    .Y(\soc/cpu/_00209_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_08596_  (.A1(\soc/cpu/_03887_ ),
    .A2(\soc/cpu/_03888_ ),
    .B1(\soc/cpu/_03886_ ),
    .Y(\soc/cpu/_03901_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08597_  (.A(\soc/cpu/decoded_imm[29] ),
    .B(\soc/cpu/reg_pc[29] ),
    .Y(\soc/cpu/_03902_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08598_  (.A(\soc/cpu/decoded_imm[29] ),
    .B(\soc/cpu/reg_pc[29] ),
    .Y(\soc/cpu/_03903_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_08599_  (.A(\soc/cpu/_03902_ ),
    .B_N(\soc/cpu/_03903_ ),
    .Y(\soc/cpu/_03904_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08600_  (.A(\soc/cpu/_03901_ ),
    .B(\soc/cpu/_03904_ ),
    .Y(\soc/cpu/_03905_ ));
 sky130_fd_sc_hd__a21boi_4 \soc/cpu/_08601_  (.A1(\soc/mem_rdata[29] ),
    .A2(net157),
    .B1_N(\soc/cpu/_03577_ ),
    .Y(\soc/cpu/_03906_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08602_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[29] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03907_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08603_  (.A1(\soc/cpu/irq_mask[29] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[29] ),
    .C1(\soc/cpu/_00872_ ),
    .Y(\soc/cpu/_03908_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08604_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[61] ),
    .B1(\soc/cpu/count_instr[29] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[61] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03909_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08605_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03909_ ),
    .Y(\soc/cpu/_03910_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08606_  (.A1(\soc/cpu/count_cycle[29] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03910_ ),
    .Y(\soc/cpu/_03911_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08607_  (.A1(\soc/cpu/_03907_ ),
    .A2(\soc/cpu/_03908_ ),
    .B1(\soc/cpu/_03911_ ),
    .Y(\soc/cpu/_03912_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08608_  (.A1(\soc/cpu/cpu_state[4] ),
    .A2(\soc/cpu/pcpi_rs1 [29]),
    .B1(\soc/cpu/_03328_ ),
    .B2(\soc/cpu/irq_pending[29] ),
    .C1(net414),
    .C2(\soc/cpu/_03912_ ),
    .Y(\soc/cpu/_03913_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08609_  (.A1(net53),
    .A2(\soc/cpu/_03906_ ),
    .B1(\soc/cpu/_03913_ ),
    .Y(\soc/cpu/_03914_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08610_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03905_ ),
    .B1(\soc/cpu/_03914_ ),
    .Y(\soc/cpu/_03915_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08611_  (.A(net131),
    .B(\soc/cpu/_03915_ ),
    .Y(\soc/cpu/_00210_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08612_  (.A(\soc/cpu/decoded_imm[30] ),
    .B(\soc/cpu/reg_pc[30] ),
    .X(\soc/cpu/_03916_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08613_  (.A(\soc/cpu/decoded_imm[30] ),
    .B(\soc/cpu/reg_pc[30] ),
    .Y(\soc/cpu/_03917_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08614_  (.A1(\soc/cpu/_03901_ ),
    .A2(\soc/cpu/_03903_ ),
    .B1(\soc/cpu/_03902_ ),
    .Y(\soc/cpu/_03918_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_08615_  (.A1(\soc/cpu/_03916_ ),
    .A2(\soc/cpu/_03917_ ),
    .B1_N(\soc/cpu/_03918_ ),
    .Y(\soc/cpu/_03919_ ));
 sky130_fd_sc_hd__a2111o_1 \soc/cpu/_08616_  (.A1(\soc/cpu/_03901_ ),
    .A2(\soc/cpu/_03903_ ),
    .B1(\soc/cpu/_03916_ ),
    .C1(\soc/cpu/_03917_ ),
    .D1(\soc/cpu/_03902_ ),
    .X(\soc/cpu/_03920_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08617_  (.A(\soc/mem_rdata[30] ),
    .B(net157),
    .Y(\soc/cpu/_03921_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08618_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03921_ ),
    .B1(net54),
    .Y(\soc/cpu/_03922_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08619_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[62] ),
    .B1(\soc/cpu/count_instr[30] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[62] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03923_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08620_  (.A1(\soc/cpu/count_cycle[30] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(net413),
    .Y(\soc/cpu/_03924_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/_08621_  (.A1(\soc/cpu/irq_mask[30] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[30] ),
    .C1(net160),
    .X(\soc/cpu/_03925_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08622_  (.A1(\soc/cpu/instr_retirq ),
    .A2(\soc/cpu/cpuregs_rdata1[30] ),
    .A3(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_03925_ ),
    .Y(\soc/cpu/_03926_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_08623_  (.A1(\soc/cpu/_03414_ ),
    .A2(\soc/cpu/_03923_ ),
    .B1(\soc/cpu/_03924_ ),
    .C1(\soc/cpu/_03926_ ),
    .Y(\soc/cpu/_03927_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08624_  (.A1(\soc/cpu/irq_pending[30] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03927_ ),
    .Y(\soc/cpu/_03928_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08625_  (.A(\soc/cpu/_02704_ ),
    .B(\soc/cpu/_03928_ ),
    .Y(\soc/cpu/_03929_ ));
 sky130_fd_sc_hd__a311oi_1 \soc/cpu/_08626_  (.A1(\soc/cpu/cpu_state[3] ),
    .A2(\soc/cpu/_03919_ ),
    .A3(\soc/cpu/_03920_ ),
    .B1(\soc/cpu/_03922_ ),
    .C1(\soc/cpu/_03929_ ),
    .Y(\soc/cpu/_03930_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08627_  (.A(net131),
    .B(\soc/cpu/_03930_ ),
    .Y(\soc/cpu/_00211_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08628_  (.A(\soc/cpu/decoded_imm[30] ),
    .B(\soc/cpu/reg_pc[30] ),
    .Y(\soc/cpu/_03931_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08629_  (.A(\soc/cpu/decoded_imm[31] ),
    .B(\soc/cpu/reg_pc[31] ),
    .Y(\soc/cpu/_03932_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08630_  (.A(\soc/cpu/_03931_ ),
    .B(\soc/cpu/_03920_ ),
    .C(\soc/cpu/_03932_ ),
    .Y(\soc/cpu/_03933_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_08631_  (.A1(\soc/cpu/_03931_ ),
    .A2(\soc/cpu/_03920_ ),
    .B1(\soc/cpu/_03932_ ),
    .X(\soc/cpu/_03934_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08632_  (.A(\soc/cpu/cpu_state[3] ),
    .B(\soc/cpu/_03933_ ),
    .C(\soc/cpu/_03934_ ),
    .Y(\soc/cpu/_03935_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08633_  (.A(\soc/cpu/cpu_state[4] ),
    .B(\soc/cpu/pcpi_rs1 [31]),
    .Y(\soc/cpu/_03936_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08634_  (.A(\soc/cpu/instr_retirq ),
    .B(\soc/cpu/cpuregs_rdata1[31] ),
    .C(\soc/cpu/_02696_ ),
    .Y(\soc/cpu/_03937_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08635_  (.A1(\soc/cpu/irq_mask[31] ),
    .A2(\soc/cpu/instr_maskirq ),
    .B1(\soc/cpu/instr_timer ),
    .B2(\soc/cpu/timer[31] ),
    .C1(\soc/cpu/_00872_ ),
    .Y(\soc/cpu/_03938_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/cpu/_08636_  (.A1(\soc/cpu/instr_rdinstrh ),
    .A2(\soc/cpu/count_instr[63] ),
    .B1(\soc/cpu/count_instr[31] ),
    .B2(\soc/cpu/instr_rdinstr ),
    .C1(\soc/cpu/count_cycle[63] ),
    .C2(\soc/cpu/instr_rdcycleh ),
    .Y(\soc/cpu/_03939_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08637_  (.A(\soc/cpu/_03414_ ),
    .B(\soc/cpu/_03939_ ),
    .Y(\soc/cpu/_03940_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/_08638_  (.A1(\soc/cpu/count_cycle[31] ),
    .A2(\soc/cpu/_00945_ ),
    .B1(\soc/cpu/_03940_ ),
    .Y(\soc/cpu/_03941_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08639_  (.A1(\soc/cpu/_03937_ ),
    .A2(\soc/cpu/_03938_ ),
    .B1(\soc/cpu/_03941_ ),
    .Y(\soc/cpu/_03942_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08640_  (.A(\soc/mem_rdata[31] ),
    .B(net157),
    .Y(\soc/cpu/_03943_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08641_  (.A1(\soc/cpu/_03577_ ),
    .A2(\soc/cpu/_03943_ ),
    .B1(net54),
    .Y(\soc/cpu/_03944_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08642_  (.A1(\soc/cpu/irq_pending[31] ),
    .A2(\soc/cpu/_03328_ ),
    .B1(\soc/cpu/_03942_ ),
    .B2(net414),
    .C1(\soc/cpu/_03944_ ),
    .Y(\soc/cpu/_03945_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08643_  (.A1(\soc/cpu/_03935_ ),
    .A2(\soc/cpu/_03936_ ),
    .A3(\soc/cpu/_03945_ ),
    .B1(net131),
    .Y(\soc/cpu/_00212_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_08644_  (.A(net413),
    .B(\soc/cpu/instr_maskirq ),
    .Y(\soc/cpu/_03946_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08647_  (.A1(\soc/cpu/irq_mask[0] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03949_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08648_  (.A1(\soc/cpu/_02916_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03949_ ),
    .Y(\soc/cpu/_00213_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08650_  (.A1(\soc/cpu/irq_mask[1] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03951_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08651_  (.A1(\soc/cpu/_02935_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03951_ ),
    .Y(\soc/cpu/_00214_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08652_  (.A1(\soc/cpu/irq_mask[2] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03952_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08653_  (.A1(\soc/cpu/_02945_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03952_ ),
    .Y(\soc/cpu/_00215_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08654_  (.A1(\soc/cpu/irq_mask[3] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03953_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08655_  (.A1(\soc/cpu/_02961_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03953_ ),
    .Y(\soc/cpu/_00216_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08656_  (.A1(\soc/cpu/irq_mask[4] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03954_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08657_  (.A1(\soc/cpu/_02980_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03954_ ),
    .Y(\soc/cpu/_00217_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08658_  (.A1(\soc/cpu/irq_mask[5] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03955_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08659_  (.A1(\soc/cpu/_02987_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03955_ ),
    .Y(\soc/cpu/_00218_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08660_  (.A1(\soc/cpu/irq_mask[6] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net132),
    .Y(\soc/cpu/_03956_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08661_  (.A1(\soc/cpu/_03008_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03956_ ),
    .Y(\soc/cpu/_00219_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08662_  (.A1(\soc/cpu/irq_mask[7] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net132),
    .Y(\soc/cpu/_03957_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08663_  (.A1(\soc/cpu/_03021_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03957_ ),
    .Y(\soc/cpu/_00220_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08665_  (.A1(\soc/cpu/irq_mask[8] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03959_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08666_  (.A1(\soc/cpu/_03033_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03959_ ),
    .Y(\soc/cpu/_00221_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08667_  (.A1(\soc/cpu/irq_mask[9] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03960_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08668_  (.A1(\soc/cpu/_03045_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03960_ ),
    .Y(\soc/cpu/_00222_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08670_  (.A1(\soc/cpu/irq_mask[10] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03962_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08671_  (.A1(\soc/cpu/_03057_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03962_ ),
    .Y(\soc/cpu/_00223_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08673_  (.A1(\soc/cpu/irq_mask[11] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03964_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08674_  (.A1(\soc/cpu/_03068_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03964_ ),
    .Y(\soc/cpu/_00224_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08675_  (.A1(\soc/cpu/irq_mask[12] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03965_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08676_  (.A1(\soc/cpu/_03076_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03965_ ),
    .Y(\soc/cpu/_00225_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08677_  (.A1(\soc/cpu/irq_mask[13] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03966_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08678_  (.A1(\soc/cpu/_03090_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03966_ ),
    .Y(\soc/cpu/_00226_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08679_  (.A1(\soc/cpu/irq_mask[14] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03967_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08680_  (.A1(\soc/cpu/_03102_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03967_ ),
    .Y(\soc/cpu/_00227_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08681_  (.A1(\soc/cpu/irq_mask[15] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03968_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08682_  (.A1(\soc/cpu/_03116_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03968_ ),
    .Y(\soc/cpu/_00228_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08683_  (.A1(\soc/cpu/irq_mask[16] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(net131),
    .Y(\soc/cpu/_03969_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08684_  (.A1(\soc/cpu/_03126_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03969_ ),
    .Y(\soc/cpu/_00229_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08685_  (.A1(\soc/cpu/irq_mask[17] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03970_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08686_  (.A1(\soc/cpu/_03136_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03970_ ),
    .Y(\soc/cpu/_00230_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08688_  (.A1(\soc/cpu/irq_mask[18] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03972_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08689_  (.A1(\soc/cpu/_03148_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03972_ ),
    .Y(\soc/cpu/_00231_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08690_  (.A1(\soc/cpu/irq_mask[19] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03973_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08691_  (.A1(\soc/cpu/_03157_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03973_ ),
    .Y(\soc/cpu/_00232_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08693_  (.A1(\soc/cpu/irq_mask[20] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03975_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08694_  (.A1(\soc/cpu/_03170_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03975_ ),
    .Y(\soc/cpu/_00233_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08696_  (.A1(\soc/cpu/irq_mask[21] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03977_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08697_  (.A1(\soc/cpu/_03180_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03977_ ),
    .Y(\soc/cpu/_00234_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08698_  (.A1(\soc/cpu/irq_mask[22] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03978_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08699_  (.A1(\soc/cpu/_03191_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03978_ ),
    .Y(\soc/cpu/_00235_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08700_  (.A1(\soc/cpu/irq_mask[23] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03979_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08701_  (.A1(\soc/cpu/_03200_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03979_ ),
    .Y(\soc/cpu/_00236_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08702_  (.A1(\soc/cpu/irq_mask[24] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03980_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08703_  (.A1(\soc/cpu/_03211_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03980_ ),
    .Y(\soc/cpu/_00237_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08704_  (.A1(\soc/cpu/irq_mask[25] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03981_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08705_  (.A1(\soc/cpu/_03223_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03981_ ),
    .Y(\soc/cpu/_00238_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08706_  (.A1(\soc/cpu/irq_mask[26] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03982_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08707_  (.A1(\soc/cpu/_03232_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03982_ ),
    .Y(\soc/cpu/_00239_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08708_  (.A1(\soc/cpu/irq_mask[27] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03983_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08709_  (.A1(\soc/cpu/_03243_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03983_ ),
    .Y(\soc/cpu/_00240_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08710_  (.A1(\soc/cpu/irq_mask[28] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03984_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08711_  (.A1(\soc/cpu/_03255_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03984_ ),
    .Y(\soc/cpu/_00241_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08712_  (.A1(\soc/cpu/irq_mask[29] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03985_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08713_  (.A1(\soc/cpu/_03267_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03985_ ),
    .Y(\soc/cpu/_00242_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08714_  (.A1(\soc/cpu/irq_mask[30] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03986_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08715_  (.A1(\soc/cpu/_03277_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03986_ ),
    .Y(\soc/cpu/_00243_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08717_  (.A1(\soc/cpu/irq_mask[31] ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_03988_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08718_  (.A1(\soc/cpu/_02698_ ),
    .A2(\soc/cpu/_03946_ ),
    .B1(\soc/cpu/_03988_ ),
    .Y(\soc/cpu/_00244_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_08719_  (.A(net413),
    .SLEEP(\soc/cpu/cpu_state[1] ),
    .X(\soc/cpu/_03989_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08720_  (.A1(\soc/cpu/irq_state[0] ),
    .A2(\soc/cpu/cpu_state[1] ),
    .B1(\soc/cpu/_03989_ ),
    .Y(\soc/cpu/_03990_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08721_  (.A1(\soc/cpu/_03397_ ),
    .A2(\soc/cpu/_03990_ ),
    .B1(\soc/cpu/irq_active ),
    .Y(\soc/cpu/_03991_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_08722_  (.A1(net413),
    .A2(\soc/cpu/_03408_ ),
    .B1(\soc/cpu/_03991_ ),
    .X(\soc/cpu/_03992_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08723_  (.A(net132),
    .B(\soc/cpu/_03992_ ),
    .Y(\soc/cpu/_00245_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_08724_  (.A(\soc/cpu/decoder_trigger ),
    .B(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_03993_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_08725_  (.A(\soc/cpu/cpu_state[1] ),
    .B(\soc/cpu/_03289_ ),
    .Y(\soc/cpu/_03994_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/_08726_  (.A(\soc/cpu/_03993_ ),
    .B(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_03995_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/_08727_  (.A0(\soc/cpu/irq_delay ),
    .A1(\soc/cpu/irq_active ),
    .S(\soc/cpu/_03995_ ),
    .Y(\soc/cpu/_03996_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08728_  (.A(net132),
    .B(\soc/cpu/_03996_ ),
    .Y(\soc/cpu/_00246_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08729_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/count_cycle[0] ),
    .Y(\soc/cpu/_00280_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08730_  (.A1(\soc/cpu/count_cycle[0] ),
    .A2(\soc/cpu/count_cycle[1] ),
    .B1(_074_),
    .Y(\soc/cpu/_03997_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08731_  (.A1(\soc/cpu/count_cycle[0] ),
    .A2(\soc/cpu/count_cycle[1] ),
    .B1(\soc/cpu/_03997_ ),
    .Y(\soc/cpu/_00281_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08732_  (.A(\soc/cpu/count_cycle[0] ),
    .B(\soc/cpu/count_cycle[1] ),
    .C(\soc/cpu/count_cycle[2] ),
    .X(\soc/cpu/_03998_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08733_  (.A1(\soc/cpu/count_cycle[0] ),
    .A2(\soc/cpu/count_cycle[1] ),
    .B1(\soc/cpu/count_cycle[2] ),
    .Y(\soc/cpu/_03999_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08734_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_03998_ ),
    .C(\soc/cpu/_03999_ ),
    .Y(\soc/cpu/_00282_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08735_  (.A(\soc/cpu/count_cycle[0] ),
    .B(\soc/cpu/count_cycle[1] ),
    .C(\soc/cpu/count_cycle[2] ),
    .D(\soc/cpu/count_cycle[3] ),
    .X(\soc/cpu/_04000_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08736_  (.A1(\soc/cpu/count_cycle[3] ),
    .A2(\soc/cpu/_03998_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04001_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08737_  (.A(\soc/cpu/_04000_ ),
    .B(\soc/cpu/_04001_ ),
    .Y(\soc/cpu/_00283_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08738_  (.A(\soc/cpu/count_cycle[4] ),
    .B(\soc/cpu/_04000_ ),
    .X(\soc/cpu/_04002_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08739_  (.A1(\soc/cpu/count_cycle[4] ),
    .A2(\soc/cpu/_04000_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04003_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08740_  (.A(\soc/cpu/_04002_ ),
    .B(\soc/cpu/_04003_ ),
    .Y(\soc/cpu/_00284_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08741_  (.A(\soc/cpu/count_cycle[4] ),
    .B(\soc/cpu/count_cycle[5] ),
    .C(\soc/cpu/_04000_ ),
    .X(\soc/cpu/_04004_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08742_  (.A1(\soc/cpu/count_cycle[5] ),
    .A2(\soc/cpu/_04002_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04005_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08743_  (.A(\soc/cpu/_04004_ ),
    .B(\soc/cpu/_04005_ ),
    .Y(\soc/cpu/_00285_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08744_  (.A1(\soc/cpu/count_cycle[6] ),
    .A2(\soc/cpu/_04004_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04006_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08745_  (.A1(\soc/cpu/count_cycle[6] ),
    .A2(\soc/cpu/_04004_ ),
    .B1(\soc/cpu/_04006_ ),
    .Y(\soc/cpu/_00286_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08746_  (.A(\soc/cpu/count_cycle[6] ),
    .B(\soc/cpu/count_cycle[7] ),
    .C(\soc/cpu/_04004_ ),
    .X(\soc/cpu/_04007_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08747_  (.A1(\soc/cpu/count_cycle[6] ),
    .A2(\soc/cpu/_04004_ ),
    .B1(\soc/cpu/count_cycle[7] ),
    .Y(\soc/cpu/_04008_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08748_  (.A(net132),
    .B(\soc/cpu/_04007_ ),
    .C(\soc/cpu/_04008_ ),
    .Y(\soc/cpu/_00287_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08749_  (.A(\soc/cpu/count_cycle[6] ),
    .B(\soc/cpu/count_cycle[7] ),
    .C(\soc/cpu/count_cycle[8] ),
    .D(\soc/cpu/_04004_ ),
    .X(\soc/cpu/_04009_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08750_  (.A1(\soc/cpu/count_cycle[8] ),
    .A2(\soc/cpu/_04007_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04010_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08751_  (.A(\soc/cpu/_04009_ ),
    .B(\soc/cpu/_04010_ ),
    .Y(\soc/cpu/_00288_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08752_  (.A(\soc/cpu/count_cycle[9] ),
    .B(\soc/cpu/_04009_ ),
    .X(\soc/cpu/_04011_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08753_  (.A1(\soc/cpu/count_cycle[9] ),
    .A2(\soc/cpu/_04009_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04012_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08754_  (.A(\soc/cpu/_04011_ ),
    .B(\soc/cpu/_04012_ ),
    .Y(\soc/cpu/_00289_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08755_  (.A(\soc/cpu/count_cycle[9] ),
    .B(\soc/cpu/count_cycle[10] ),
    .C(\soc/cpu/_04009_ ),
    .X(\soc/cpu/_04013_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08756_  (.A1(\soc/cpu/count_cycle[10] ),
    .A2(\soc/cpu/_04011_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04014_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08757_  (.A(\soc/cpu/_04013_ ),
    .B(\soc/cpu/_04014_ ),
    .Y(\soc/cpu/_00290_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08758_  (.A(\soc/cpu/count_cycle[9] ),
    .B(\soc/cpu/count_cycle[10] ),
    .C(\soc/cpu/count_cycle[11] ),
    .D(\soc/cpu/_04009_ ),
    .X(\soc/cpu/_04015_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08759_  (.A1(\soc/cpu/count_cycle[11] ),
    .A2(\soc/cpu/_04013_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04016_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08760_  (.A(\soc/cpu/_04015_ ),
    .B(\soc/cpu/_04016_ ),
    .Y(\soc/cpu/_00291_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08761_  (.A1(\soc/cpu/count_cycle[12] ),
    .A2(\soc/cpu/_04015_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04017_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08762_  (.A1(\soc/cpu/count_cycle[12] ),
    .A2(\soc/cpu/_04015_ ),
    .B1(\soc/cpu/_04017_ ),
    .Y(\soc/cpu/_00292_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08763_  (.A(\soc/cpu/count_cycle[12] ),
    .B(\soc/cpu/count_cycle[13] ),
    .C(\soc/cpu/_04015_ ),
    .X(\soc/cpu/_04018_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08764_  (.A1(\soc/cpu/count_cycle[12] ),
    .A2(\soc/cpu/_04015_ ),
    .B1(\soc/cpu/count_cycle[13] ),
    .Y(\soc/cpu/_04019_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08765_  (.A(net132),
    .B(\soc/cpu/_04018_ ),
    .C(\soc/cpu/_04019_ ),
    .Y(\soc/cpu/_00293_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08766_  (.A(\soc/cpu/count_cycle[12] ),
    .B(\soc/cpu/count_cycle[13] ),
    .C(\soc/cpu/count_cycle[14] ),
    .D(\soc/cpu/_04015_ ),
    .X(\soc/cpu/_04020_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08767_  (.A1(\soc/cpu/count_cycle[14] ),
    .A2(\soc/cpu/_04018_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04021_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08768_  (.A(\soc/cpu/_04020_ ),
    .B(\soc/cpu/_04021_ ),
    .Y(\soc/cpu/_00294_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08769_  (.A(\soc/cpu/count_cycle[15] ),
    .B(\soc/cpu/_04020_ ),
    .X(\soc/cpu/_04022_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08770_  (.A1(\soc/cpu/count_cycle[15] ),
    .A2(\soc/cpu/_04020_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04023_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08771_  (.A(\soc/cpu/_04022_ ),
    .B(\soc/cpu/_04023_ ),
    .Y(\soc/cpu/_00295_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08772_  (.A(\soc/cpu/count_cycle[15] ),
    .B(\soc/cpu/count_cycle[16] ),
    .C(\soc/cpu/_04020_ ),
    .X(\soc/cpu/_04024_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08774_  (.A1(\soc/cpu/count_cycle[16] ),
    .A2(\soc/cpu/_04022_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04026_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08775_  (.A(\soc/cpu/_04024_ ),
    .B(\soc/cpu/_04026_ ),
    .Y(\soc/cpu/_00296_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08776_  (.A(\soc/cpu/count_cycle[15] ),
    .B(\soc/cpu/count_cycle[16] ),
    .C(\soc/cpu/count_cycle[17] ),
    .D(\soc/cpu/_04020_ ),
    .X(\soc/cpu/_04027_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08777_  (.A1(\soc/cpu/count_cycle[17] ),
    .A2(\soc/cpu/_04024_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04028_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08778_  (.A(\soc/cpu/_04027_ ),
    .B(\soc/cpu/_04028_ ),
    .Y(\soc/cpu/_00297_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08780_  (.A1(\soc/cpu/count_cycle[18] ),
    .A2(\soc/cpu/_04027_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04030_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08781_  (.A1(\soc/cpu/count_cycle[18] ),
    .A2(\soc/cpu/_04027_ ),
    .B1(\soc/cpu/_04030_ ),
    .Y(\soc/cpu/_00298_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08782_  (.A(\soc/cpu/count_cycle[18] ),
    .B(\soc/cpu/count_cycle[19] ),
    .C(\soc/cpu/_04027_ ),
    .X(\soc/cpu/_04031_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08783_  (.A1(\soc/cpu/count_cycle[18] ),
    .A2(\soc/cpu/_04027_ ),
    .B1(\soc/cpu/count_cycle[19] ),
    .Y(\soc/cpu/_04032_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08784_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04031_ ),
    .C(\soc/cpu/_04032_ ),
    .Y(\soc/cpu/_00299_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08785_  (.A(\soc/cpu/count_cycle[18] ),
    .B(\soc/cpu/count_cycle[19] ),
    .C(\soc/cpu/count_cycle[20] ),
    .D(\soc/cpu/_04027_ ),
    .X(\soc/cpu/_04033_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08786_  (.A1(\soc/cpu/count_cycle[20] ),
    .A2(\soc/cpu/_04031_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04034_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08787_  (.A(\soc/cpu/_04033_ ),
    .B(\soc/cpu/_04034_ ),
    .Y(\soc/cpu/_00300_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08788_  (.A(\soc/cpu/count_cycle[21] ),
    .B(\soc/cpu/_04033_ ),
    .X(\soc/cpu/_04035_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08789_  (.A(\soc/cpu/count_cycle[21] ),
    .B(\soc/cpu/_04033_ ),
    .Y(\soc/cpu/_04036_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08790_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04035_ ),
    .C(\soc/cpu/_04036_ ),
    .Y(\soc/cpu/_00301_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08791_  (.A(\soc/cpu/count_cycle[21] ),
    .B(\soc/cpu/count_cycle[22] ),
    .C(\soc/cpu/_04033_ ),
    .X(\soc/cpu/_04037_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08792_  (.A1(\soc/cpu/count_cycle[22] ),
    .A2(\soc/cpu/_04035_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04038_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08793_  (.A(\soc/cpu/_04037_ ),
    .B(\soc/cpu/_04038_ ),
    .Y(\soc/cpu/_00302_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08794_  (.A(\soc/cpu/count_cycle[21] ),
    .B(\soc/cpu/count_cycle[22] ),
    .C(\soc/cpu/count_cycle[23] ),
    .D(\soc/cpu/_04033_ ),
    .X(\soc/cpu/_04039_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08795_  (.A1(\soc/cpu/count_cycle[23] ),
    .A2(\soc/cpu/_04037_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04040_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08796_  (.A(\soc/cpu/_04039_ ),
    .B(\soc/cpu/_04040_ ),
    .Y(\soc/cpu/_00303_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08797_  (.A1(\soc/cpu/count_cycle[24] ),
    .A2(\soc/cpu/_04039_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04041_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08798_  (.A1(\soc/cpu/count_cycle[24] ),
    .A2(\soc/cpu/_04039_ ),
    .B1(\soc/cpu/_04041_ ),
    .Y(\soc/cpu/_00304_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08799_  (.A(\soc/cpu/count_cycle[24] ),
    .B(\soc/cpu/count_cycle[25] ),
    .C(\soc/cpu/_04039_ ),
    .X(\soc/cpu/_04042_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08800_  (.A1(\soc/cpu/count_cycle[24] ),
    .A2(\soc/cpu/_04039_ ),
    .B1(\soc/cpu/count_cycle[25] ),
    .Y(\soc/cpu/_04043_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08801_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04042_ ),
    .C(\soc/cpu/_04043_ ),
    .Y(\soc/cpu/_00305_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08802_  (.A(\soc/cpu/count_cycle[24] ),
    .B(\soc/cpu/count_cycle[25] ),
    .C(\soc/cpu/count_cycle[26] ),
    .D(\soc/cpu/_04039_ ),
    .X(\soc/cpu/_04044_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08803_  (.A1(\soc/cpu/count_cycle[26] ),
    .A2(\soc/cpu/_04042_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04045_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08804_  (.A(\soc/cpu/_04044_ ),
    .B(\soc/cpu/_04045_ ),
    .Y(\soc/cpu/_00306_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08805_  (.A(\soc/cpu/count_cycle[27] ),
    .B(\soc/cpu/_04044_ ),
    .X(\soc/cpu/_04046_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08806_  (.A(\soc/cpu/count_cycle[27] ),
    .B(\soc/cpu/_04044_ ),
    .Y(\soc/cpu/_04047_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08807_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04046_ ),
    .C(\soc/cpu/_04047_ ),
    .Y(\soc/cpu/_00307_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08808_  (.A(\soc/cpu/count_cycle[27] ),
    .B(\soc/cpu/count_cycle[28] ),
    .C(\soc/cpu/_04044_ ),
    .X(\soc/cpu/_04048_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08809_  (.A1(\soc/cpu/count_cycle[28] ),
    .A2(\soc/cpu/_04046_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04049_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08810_  (.A(\soc/cpu/_04048_ ),
    .B(\soc/cpu/_04049_ ),
    .Y(\soc/cpu/_00308_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08811_  (.A(\soc/cpu/count_cycle[27] ),
    .B(\soc/cpu/count_cycle[28] ),
    .C(\soc/cpu/count_cycle[29] ),
    .D(\soc/cpu/_04044_ ),
    .X(\soc/cpu/_04050_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08812_  (.A1(\soc/cpu/count_cycle[29] ),
    .A2(\soc/cpu/_04048_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04051_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08813_  (.A(\soc/cpu/_04050_ ),
    .B(\soc/cpu/_04051_ ),
    .Y(\soc/cpu/_00309_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08814_  (.A1(\soc/cpu/count_cycle[30] ),
    .A2(\soc/cpu/_04050_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04052_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08815_  (.A1(\soc/cpu/count_cycle[30] ),
    .A2(\soc/cpu/_04050_ ),
    .B1(\soc/cpu/_04052_ ),
    .Y(\soc/cpu/_00310_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08816_  (.A(\soc/cpu/count_cycle[30] ),
    .B(\soc/cpu/count_cycle[31] ),
    .C(\soc/cpu/_04050_ ),
    .X(\soc/cpu/_04053_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08817_  (.A1(\soc/cpu/count_cycle[30] ),
    .A2(\soc/cpu/_04050_ ),
    .B1(\soc/cpu/count_cycle[31] ),
    .Y(\soc/cpu/_04054_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08818_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04053_ ),
    .C(\soc/cpu/_04054_ ),
    .Y(\soc/cpu/_00311_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08819_  (.A(\soc/cpu/count_cycle[32] ),
    .B(\soc/cpu/count_cycle[30] ),
    .C(\soc/cpu/count_cycle[31] ),
    .D(\soc/cpu/_04050_ ),
    .X(\soc/cpu/_04055_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08820_  (.A1(\soc/cpu/count_cycle[32] ),
    .A2(\soc/cpu/_04053_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04056_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08821_  (.A(\soc/cpu/_04055_ ),
    .B(\soc/cpu/_04056_ ),
    .Y(\soc/cpu/_00312_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08822_  (.A(\soc/cpu/count_cycle[33] ),
    .B(\soc/cpu/_04055_ ),
    .X(\soc/cpu/_04057_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08823_  (.A(\soc/cpu/count_cycle[33] ),
    .B(\soc/cpu/_04055_ ),
    .Y(\soc/cpu/_04058_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08824_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04057_ ),
    .C(\soc/cpu/_04058_ ),
    .Y(\soc/cpu/_00313_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08825_  (.A(\soc/cpu/count_cycle[33] ),
    .B(\soc/cpu/count_cycle[34] ),
    .C(\soc/cpu/_04055_ ),
    .X(\soc/cpu/_04059_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08826_  (.A1(\soc/cpu/count_cycle[34] ),
    .A2(\soc/cpu/_04057_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04060_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08827_  (.A(\soc/cpu/_04059_ ),
    .B(\soc/cpu/_04060_ ),
    .Y(\soc/cpu/_00314_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08828_  (.A(\soc/cpu/count_cycle[33] ),
    .B(\soc/cpu/count_cycle[34] ),
    .C(\soc/cpu/count_cycle[35] ),
    .D(\soc/cpu/_04055_ ),
    .X(\soc/cpu/_04061_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08830_  (.A1(\soc/cpu/count_cycle[35] ),
    .A2(\soc/cpu/_04059_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04063_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08831_  (.A(\soc/cpu/_04061_ ),
    .B(\soc/cpu/_04063_ ),
    .Y(\soc/cpu/_00315_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08832_  (.A1(\soc/cpu/count_cycle[36] ),
    .A2(\soc/cpu/_04061_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04064_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08833_  (.A1(\soc/cpu/count_cycle[36] ),
    .A2(\soc/cpu/_04061_ ),
    .B1(\soc/cpu/_04064_ ),
    .Y(\soc/cpu/_00316_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08835_  (.A(\soc/cpu/count_cycle[36] ),
    .B(\soc/cpu/count_cycle[37] ),
    .C(\soc/cpu/_04061_ ),
    .X(\soc/cpu/_04066_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08836_  (.A1(\soc/cpu/count_cycle[36] ),
    .A2(\soc/cpu/_04061_ ),
    .B1(\soc/cpu/count_cycle[37] ),
    .Y(\soc/cpu/_04067_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08837_  (.A(net132),
    .B(\soc/cpu/_04066_ ),
    .C(\soc/cpu/_04067_ ),
    .Y(\soc/cpu/_00317_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08838_  (.A(\soc/cpu/count_cycle[36] ),
    .B(\soc/cpu/count_cycle[37] ),
    .C(\soc/cpu/count_cycle[38] ),
    .D(\soc/cpu/_04061_ ),
    .X(\soc/cpu/_04068_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08839_  (.A1(\soc/cpu/count_cycle[38] ),
    .A2(\soc/cpu/_04066_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04069_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08840_  (.A(\soc/cpu/_04068_ ),
    .B(\soc/cpu/_04069_ ),
    .Y(\soc/cpu/_00318_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08841_  (.A(\soc/cpu/count_cycle[39] ),
    .B(\soc/cpu/_04068_ ),
    .X(\soc/cpu/_04070_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08842_  (.A1(\soc/cpu/count_cycle[39] ),
    .A2(\soc/cpu/_04068_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04071_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08843_  (.A(\soc/cpu/_04070_ ),
    .B(\soc/cpu/_04071_ ),
    .Y(\soc/cpu/_00319_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08844_  (.A(\soc/cpu/count_cycle[39] ),
    .B(\soc/cpu/count_cycle[40] ),
    .C(\soc/cpu/_04068_ ),
    .X(\soc/cpu/_04072_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08845_  (.A1(\soc/cpu/count_cycle[40] ),
    .A2(\soc/cpu/_04070_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04073_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08846_  (.A(\soc/cpu/_04072_ ),
    .B(\soc/cpu/_04073_ ),
    .Y(\soc/cpu/_00320_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08847_  (.A(\soc/cpu/count_cycle[39] ),
    .B(\soc/cpu/count_cycle[40] ),
    .C(\soc/cpu/count_cycle[41] ),
    .D(\soc/cpu/_04068_ ),
    .X(\soc/cpu/_04074_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08848_  (.A1(\soc/cpu/count_cycle[41] ),
    .A2(\soc/cpu/_04072_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04075_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08849_  (.A(\soc/cpu/_04074_ ),
    .B(\soc/cpu/_04075_ ),
    .Y(\soc/cpu/_00321_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08850_  (.A1(\soc/cpu/count_cycle[42] ),
    .A2(\soc/cpu/_04074_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04076_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08851_  (.A1(\soc/cpu/count_cycle[42] ),
    .A2(\soc/cpu/_04074_ ),
    .B1(\soc/cpu/_04076_ ),
    .Y(\soc/cpu/_00322_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08852_  (.A(\soc/cpu/count_cycle[42] ),
    .B(net789),
    .C(\soc/cpu/_04074_ ),
    .X(\soc/cpu/_04077_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08853_  (.A1(\soc/cpu/count_cycle[42] ),
    .A2(\soc/cpu/_04074_ ),
    .B1(\soc/cpu/count_cycle[43] ),
    .Y(\soc/cpu/_04078_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08854_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04077_ ),
    .C(\soc/cpu/_04078_ ),
    .Y(\soc/cpu/_00323_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08855_  (.A(net795),
    .B(net789),
    .C(\soc/cpu/count_cycle[44] ),
    .D(\soc/cpu/_04074_ ),
    .X(\soc/cpu/_04079_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08856_  (.A1(\soc/cpu/count_cycle[44] ),
    .A2(net790),
    .B1(_074_),
    .Y(\soc/cpu/_04080_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08857_  (.A(\soc/cpu/_04079_ ),
    .B(\soc/cpu/_04080_ ),
    .Y(\soc/cpu/_00324_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08858_  (.A(\soc/cpu/count_cycle[45] ),
    .B(\soc/cpu/_04079_ ),
    .X(\soc/cpu/_04081_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08859_  (.A(\soc/cpu/count_cycle[45] ),
    .B(\soc/cpu/_04079_ ),
    .Y(\soc/cpu/_04082_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08860_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04081_ ),
    .C(\soc/cpu/_04082_ ),
    .Y(\soc/cpu/_00325_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08861_  (.A(\soc/cpu/count_cycle[45] ),
    .B(\soc/cpu/count_cycle[46] ),
    .C(\soc/cpu/_04079_ ),
    .X(\soc/cpu/_04083_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08862_  (.A1(\soc/cpu/count_cycle[46] ),
    .A2(\soc/cpu/_04081_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04084_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08863_  (.A(\soc/cpu/_04083_ ),
    .B(\soc/cpu/_04084_ ),
    .Y(\soc/cpu/_00326_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08864_  (.A(\soc/cpu/count_cycle[45] ),
    .B(\soc/cpu/count_cycle[46] ),
    .C(\soc/cpu/count_cycle[47] ),
    .D(\soc/cpu/_04079_ ),
    .X(\soc/cpu/_04085_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08865_  (.A1(\soc/cpu/count_cycle[47] ),
    .A2(\soc/cpu/_04083_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04086_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08866_  (.A(\soc/cpu/_04085_ ),
    .B(\soc/cpu/_04086_ ),
    .Y(\soc/cpu/_00327_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08867_  (.A1(\soc/cpu/count_cycle[48] ),
    .A2(\soc/cpu/_04085_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04087_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08868_  (.A1(\soc/cpu/count_cycle[48] ),
    .A2(\soc/cpu/_04085_ ),
    .B1(\soc/cpu/_04087_ ),
    .Y(\soc/cpu/_00328_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08869_  (.A(\soc/cpu/count_cycle[48] ),
    .B(\soc/cpu/count_cycle[49] ),
    .C(\soc/cpu/_04085_ ),
    .X(\soc/cpu/_04088_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08870_  (.A1(\soc/cpu/count_cycle[48] ),
    .A2(\soc/cpu/_04085_ ),
    .B1(\soc/cpu/count_cycle[49] ),
    .Y(\soc/cpu/_04089_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08871_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04088_ ),
    .C(\soc/cpu/_04089_ ),
    .Y(\soc/cpu/_00329_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08872_  (.A1(\soc/cpu/count_cycle[50] ),
    .A2(\soc/cpu/_04088_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04090_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08873_  (.A1(\soc/cpu/count_cycle[50] ),
    .A2(\soc/cpu/_04088_ ),
    .B1(\soc/cpu/_04090_ ),
    .Y(\soc/cpu/_00330_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08874_  (.A(\soc/cpu/count_cycle[50] ),
    .B(\soc/cpu/count_cycle[51] ),
    .C(\soc/cpu/_04088_ ),
    .X(\soc/cpu/_04091_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08875_  (.A1(\soc/cpu/count_cycle[50] ),
    .A2(\soc/cpu/_04088_ ),
    .B1(\soc/cpu/count_cycle[51] ),
    .Y(\soc/cpu/_04092_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08876_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04091_ ),
    .C(\soc/cpu/_04092_ ),
    .Y(\soc/cpu/_00331_ ));
 sky130_fd_sc_hd__and4_2 \soc/cpu/_08877_  (.A(\soc/cpu/count_cycle[50] ),
    .B(\soc/cpu/count_cycle[51] ),
    .C(\soc/cpu/count_cycle[52] ),
    .D(\soc/cpu/_04088_ ),
    .X(\soc/cpu/_04093_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08878_  (.A1(\soc/cpu/count_cycle[52] ),
    .A2(\soc/cpu/_04091_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04094_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08879_  (.A(\soc/cpu/_04093_ ),
    .B(\soc/cpu/_04094_ ),
    .Y(\soc/cpu/_00332_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08880_  (.A1(\soc/cpu/count_cycle[53] ),
    .A2(\soc/cpu/_04093_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04095_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08881_  (.A1(\soc/cpu/count_cycle[53] ),
    .A2(\soc/cpu/_04093_ ),
    .B1(\soc/cpu/_04095_ ),
    .Y(\soc/cpu/_00333_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08882_  (.A(\soc/cpu/count_cycle[53] ),
    .B(\soc/cpu/count_cycle[54] ),
    .C(\soc/cpu/_04093_ ),
    .X(\soc/cpu/_04096_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08883_  (.A1(\soc/cpu/count_cycle[53] ),
    .A2(\soc/cpu/_04093_ ),
    .B1(\soc/cpu/count_cycle[54] ),
    .Y(\soc/cpu/_04097_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08884_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04096_ ),
    .C(\soc/cpu/_04097_ ),
    .Y(\soc/cpu/_00334_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_08885_  (.A(\soc/cpu/count_cycle[53] ),
    .B(\soc/cpu/count_cycle[54] ),
    .C(\soc/cpu/count_cycle[55] ),
    .D(\soc/cpu/_04093_ ),
    .X(\soc/cpu/_04098_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08886_  (.A1(\soc/cpu/count_cycle[53] ),
    .A2(\soc/cpu/count_cycle[54] ),
    .A3(\soc/cpu/_04093_ ),
    .B1(\soc/cpu/count_cycle[55] ),
    .Y(\soc/cpu/_04099_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08887_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04098_ ),
    .C(\soc/cpu/_04099_ ),
    .Y(\soc/cpu/_00335_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08888_  (.A1(\soc/cpu/count_cycle[56] ),
    .A2(\soc/cpu/_04098_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04100_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08889_  (.A1(\soc/cpu/count_cycle[56] ),
    .A2(\soc/cpu/_04098_ ),
    .B1(\soc/cpu/_04100_ ),
    .Y(\soc/cpu/_00336_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08890_  (.A(\soc/cpu/count_cycle[56] ),
    .B(\soc/cpu/count_cycle[57] ),
    .C(\soc/cpu/_04098_ ),
    .X(\soc/cpu/_04101_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08891_  (.A1(\soc/cpu/count_cycle[56] ),
    .A2(\soc/cpu/_04098_ ),
    .B1(\soc/cpu/count_cycle[57] ),
    .Y(\soc/cpu/_04102_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08892_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04101_ ),
    .C(\soc/cpu/_04102_ ),
    .Y(\soc/cpu/_00337_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_08893_  (.A(\soc/cpu/count_cycle[58] ),
    .B(\soc/cpu/_04101_ ),
    .X(\soc/cpu/_04103_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08894_  (.A1(\soc/cpu/count_cycle[58] ),
    .A2(\soc/cpu/_04101_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04104_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08895_  (.A(\soc/cpu/_04103_ ),
    .B(\soc/cpu/_04104_ ),
    .Y(\soc/cpu/_00338_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08896_  (.A1(\soc/cpu/count_cycle[59] ),
    .A2(\soc/cpu/_04103_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04105_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08897_  (.A1(\soc/cpu/count_cycle[59] ),
    .A2(\soc/cpu/_04103_ ),
    .B1(\soc/cpu/_04105_ ),
    .Y(\soc/cpu/_00339_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08898_  (.A1(\soc/cpu/count_cycle[59] ),
    .A2(\soc/cpu/_04103_ ),
    .B1(\soc/cpu/count_cycle[60] ),
    .Y(\soc/cpu/_04106_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08899_  (.A(\soc/cpu/count_cycle[59] ),
    .B(\soc/cpu/count_cycle[60] ),
    .C(\soc/cpu/_04103_ ),
    .Y(\soc/cpu/_04107_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/cpu/_08900_  (.A(\soc/cpu/_04106_ ),
    .B(\soc/cpu/_00840_ ),
    .C_N(\soc/cpu/_04107_ ),
    .Y(\soc/cpu/_00340_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/cpu/_08901_  (.A(\soc/cpu/count_cycle[61] ),
    .SLEEP(\soc/cpu/_04107_ ),
    .X(\soc/cpu/_04108_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_08902_  (.A1(\soc/cpu/count_cycle[59] ),
    .A2(\soc/cpu/count_cycle[60] ),
    .A3(\soc/cpu/_04103_ ),
    .B1(\soc/cpu/count_cycle[61] ),
    .Y(\soc/cpu/_04109_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08903_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04108_ ),
    .C(\soc/cpu/_04109_ ),
    .Y(\soc/cpu/_00341_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08905_  (.A1(\soc/cpu/count_cycle[62] ),
    .A2(\soc/cpu/_04108_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04111_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08906_  (.A1(\soc/cpu/count_cycle[62] ),
    .A2(\soc/cpu/_04108_ ),
    .B1(\soc/cpu/_04111_ ),
    .Y(\soc/cpu/_00342_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08907_  (.A(\soc/cpu/count_cycle[62] ),
    .B(\soc/cpu/count_cycle[63] ),
    .C(\soc/cpu/_04108_ ),
    .X(\soc/cpu/_04112_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08908_  (.A1(\soc/cpu/count_cycle[62] ),
    .A2(\soc/cpu/_04108_ ),
    .B1(\soc/cpu/count_cycle[63] ),
    .Y(\soc/cpu/_04113_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_08909_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04112_ ),
    .C(\soc/cpu/_04113_ ),
    .Y(\soc/cpu/_00343_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_08910_  (.A(\soc/cpu/_00839_ ),
    .B(\soc/cpu/_03289_ ),
    .Y(\soc/cpu/_04114_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/_08912_  (.A0(\soc/cpu/irq_state[0] ),
    .A1(\soc/cpu/latched_store ),
    .S(\soc/cpu/latched_branch ),
    .Y(\soc/cpu/_04116_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08914_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02124_ ),
    .B1(\soc/cpu/_04116_ ),
    .Y(\soc/cpu/_04118_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08915_  (.A(\soc/cpu/_00708_ ),
    .B(\soc/cpu/_04118_ ),
    .Y(\soc/cpu/_04119_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08916_  (.A(\soc/cpu/_04114_ ),
    .B(\soc/cpu/_04119_ ),
    .Y(\soc/cpu/_04120_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_08917_  (.A1(\soc/cpu/latched_store ),
    .A2(\soc/cpu/latched_branch ),
    .B1(\soc/cpu/reg_next_pc[1] ),
    .X(\soc/cpu/_04121_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/_08918_  (.A1(\soc/cpu/latched_branch ),
    .A2(\soc/cpu/_02143_ ),
    .B1(\soc/cpu/_00709_ ),
    .B2(\soc/cpu/_02124_ ),
    .C1(\soc/cpu/_04121_ ),
    .Y(\soc/cpu/_04122_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_08919_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_03993_ ),
    .B1(\soc/cpu/_03403_ ),
    .Y(\soc/cpu/_04123_ ));
 sky130_fd_sc_hd__a32oi_2 \soc/cpu/_08920_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/decoded_imm_j[1] ),
    .A3(\soc/cpu/_00928_ ),
    .B1(\soc/cpu/_04123_ ),
    .B2(\soc/cpu/compressed_instr ),
    .Y(\soc/cpu/_04124_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08921_  (.A1(\soc/cpu/compressed_instr ),
    .A2(\soc/cpu/_03403_ ),
    .B1(\soc/cpu/_04119_ ),
    .Y(\soc/cpu/_04125_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/cpu/_08922_  (.A1(\soc/cpu/_04124_ ),
    .A2(\soc/cpu/_04125_ ),
    .B1_N(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04126_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08923_  (.A1(\soc/cpu/_04122_ ),
    .A2(\soc/cpu/_04124_ ),
    .B1(\soc/cpu/_04126_ ),
    .Y(\soc/cpu/_04127_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08924_  (.A1(\soc/cpu/reg_next_pc[1] ),
    .A2(\soc/cpu/_00839_ ),
    .B1(\soc/cpu/_04127_ ),
    .Y(\soc/cpu/_04128_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08925_  (.A1(\soc/cpu/_04120_ ),
    .A2(\soc/cpu/_04128_ ),
    .B1(net132),
    .Y(\soc/cpu/_00344_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_08927_  (.A(\soc/cpu/compressed_instr ),
    .B(\soc/cpu/_04122_ ),
    .C(\soc/cpu/_04123_ ),
    .X(\soc/cpu/_04130_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_08928_  (.A(\soc/cpu/_00928_ ),
    .B(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04131_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_08930_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02132_ ),
    .B1(\soc/cpu/_04116_ ),
    .B2(\soc/cpu/reg_next_pc[2] ),
    .Y(\soc/cpu/_04133_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08931_  (.A1(\soc/cpu/_04130_ ),
    .A2(\soc/cpu/_04131_ ),
    .B1(\soc/cpu/_04133_ ),
    .Y(\soc/cpu/_04134_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08932_  (.A(\soc/cpu/_02444_ ),
    .B(\soc/cpu/_04122_ ),
    .Y(\soc/cpu/_04135_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/cpu/_08933_  (.A_N(\soc/cpu/latched_branch ),
    .B(\soc/cpu/irq_state[0] ),
    .Y(\soc/cpu/_04136_ ));
 sky130_fd_sc_hd__o2111ai_4 \soc/cpu/_08934_  (.A1(\soc/cpu/_00709_ ),
    .A2(\soc/cpu/_02132_ ),
    .B1(\soc/cpu/_04136_ ),
    .C1(\soc/cpu/_01597_ ),
    .D1(\soc/cpu/decoded_imm_j[2] ),
    .Y(\soc/cpu/_04137_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_08935_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02132_ ),
    .B1(\soc/cpu/_04116_ ),
    .B2(\soc/cpu/reg_next_pc[2] ),
    .C1(\soc/cpu/decoded_imm_j[2] ),
    .Y(\soc/cpu/_04138_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_08936_  (.A(\soc/cpu/_04137_ ),
    .SLEEP(\soc/cpu/_04138_ ),
    .X(\soc/cpu/_04139_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08937_  (.A(\soc/cpu/_04135_ ),
    .B(\soc/cpu/_04139_ ),
    .Y(\soc/cpu/_04140_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08938_  (.A1(\soc/cpu/compressed_instr ),
    .A2(\soc/cpu/_04122_ ),
    .B1(\soc/cpu/_04133_ ),
    .Y(\soc/cpu/_04141_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08940_  (.A1(\soc/cpu/_03312_ ),
    .A2(\soc/cpu/_04140_ ),
    .B1(\soc/cpu/_04141_ ),
    .B2(\soc/cpu/_04123_ ),
    .C1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04143_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08941_  (.A(\soc/cpu/_00953_ ),
    .B(\soc/cpu/_04133_ ),
    .Y(\soc/cpu/_04144_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08942_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[2] ),
    .B1(\soc/cpu/_04134_ ),
    .B2(\soc/cpu/_04143_ ),
    .C1(\soc/cpu/_04144_ ),
    .Y(\soc/cpu/_04145_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08943_  (.A(net132),
    .B(\soc/cpu/_04145_ ),
    .Y(\soc/cpu/_00345_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/_08944_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02136_ ),
    .B1(\soc/cpu/_04116_ ),
    .B2(\soc/cpu/_01606_ ),
    .Y(\soc/cpu/_04146_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08945_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_00797_ ),
    .B1(\soc/cpu/_04141_ ),
    .Y(\soc/cpu/_04147_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_08946_  (.A(\soc/cpu/_00791_ ),
    .B(\soc/cpu/_04131_ ),
    .C(\soc/cpu/_04147_ ),
    .X(\soc/cpu/_04148_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08947_  (.A1(\soc/cpu/cpu_state[1] ),
    .A2(\soc/cpu/reg_next_pc[3] ),
    .B1(_074_),
    .Y(\soc/cpu/_04149_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/_08948_  (.A1(\soc/cpu/_02444_ ),
    .A2(\soc/cpu/_04122_ ),
    .A3(\soc/cpu/_04138_ ),
    .B1(\soc/cpu/_04137_ ),
    .Y(\soc/cpu/_04150_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08949_  (.A(\soc/cpu/_02454_ ),
    .B(\soc/cpu/_04146_ ),
    .Y(\soc/cpu/_04151_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08950_  (.A(\soc/cpu/_02454_ ),
    .B(\soc/cpu/_04146_ ),
    .Y(\soc/cpu/_04152_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_08951_  (.A(\soc/cpu/_04151_ ),
    .SLEEP(\soc/cpu/_04152_ ),
    .X(\soc/cpu/_04153_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08952_  (.A(\soc/cpu/_04150_ ),
    .B(\soc/cpu/_04153_ ),
    .Y(\soc/cpu/_04154_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08953_  (.A(\soc/cpu/_03312_ ),
    .B(\soc/cpu/_04154_ ),
    .Y(\soc/cpu/_04155_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/cpu/_08954_  (.A1(\soc/cpu/compressed_instr ),
    .A2(\soc/cpu/_04122_ ),
    .B1(\soc/cpu/_04133_ ),
    .C1(\soc/cpu/_04146_ ),
    .Y(\soc/cpu/_04156_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08955_  (.A(\soc/cpu/_04123_ ),
    .B(\soc/cpu/_04156_ ),
    .Y(\soc/cpu/_04157_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08957_  (.A1(\soc/cpu/_04155_ ),
    .A2(\soc/cpu/_04157_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04159_ ));
 sky130_fd_sc_hd__a311oi_1 \soc/cpu/_08958_  (.A1(\soc/cpu/cpu_state[1] ),
    .A2(\soc/cpu/_04146_ ),
    .A3(\soc/cpu/_04148_ ),
    .B1(\soc/cpu/_04149_ ),
    .C1(\soc/cpu/_04159_ ),
    .Y(\soc/cpu/_00346_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08959_  (.A1(\soc/cpu/_04150_ ),
    .A2(\soc/cpu/_04151_ ),
    .B1(\soc/cpu/_04152_ ),
    .Y(\soc/cpu/_04160_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08960_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02142_ ),
    .B1(\soc/cpu/_04116_ ),
    .Y(\soc/cpu/_04161_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08961_  (.A1(\soc/cpu/_02144_ ),
    .A2(\soc/cpu/_00709_ ),
    .B1(\soc/cpu/_04161_ ),
    .Y(\soc/cpu/_04162_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_08962_  (.A(\soc/cpu/decoded_imm_j[4] ),
    .B(\soc/cpu/_04162_ ),
    .X(\soc/cpu/_04163_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08963_  (.A(\soc/cpu/_04160_ ),
    .B(\soc/cpu/_04163_ ),
    .Y(\soc/cpu/_04164_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08964_  (.A(\soc/cpu/_04157_ ),
    .B(\soc/cpu/_04162_ ),
    .Y(\soc/cpu/_04165_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08965_  (.A1(\soc/cpu/_03312_ ),
    .A2(\soc/cpu/_04164_ ),
    .B1(\soc/cpu/_04165_ ),
    .Y(\soc/cpu/_04166_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08966_  (.A(\soc/cpu/_04156_ ),
    .B(\soc/cpu/_04162_ ),
    .Y(\soc/cpu/_04167_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/_08967_  (.A1(\soc/cpu/_04123_ ),
    .A2(\soc/cpu/_04167_ ),
    .B1(\soc/cpu/_04131_ ),
    .C1(\soc/cpu/_00791_ ),
    .X(\soc/cpu/_04168_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_08968_  (.A(\soc/cpu/cpu_state[1] ),
    .B(\soc/cpu/_04162_ ),
    .C(\soc/cpu/_04168_ ),
    .Y(\soc/cpu/_04169_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/_08969_  (.A1(\soc/cpu/cpu_state[1] ),
    .A2(\soc/cpu/_02144_ ),
    .B1(\soc/cpu/_03994_ ),
    .B2(\soc/cpu/_04166_ ),
    .C1(\soc/cpu/_04169_ ),
    .Y(\soc/cpu/_04170_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_08970_  (.A(_074_),
    .B(\soc/cpu/_04170_ ),
    .X(\soc/cpu/_00347_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08971_  (.A1(\soc/cpu/reg_next_pc[5] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04171_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08972_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02152_ ),
    .B1(\soc/cpu/_04171_ ),
    .Y(\soc/cpu/_04172_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08973_  (.A(\soc/cpu/_04167_ ),
    .B(\soc/cpu/_04172_ ),
    .Y(\soc/cpu/_04173_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08974_  (.A(\soc/cpu/_04123_ ),
    .B(\soc/cpu/_04173_ ),
    .Y(\soc/cpu/_04174_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08975_  (.A(\soc/cpu/decoded_imm_j[5] ),
    .B(\soc/cpu/_04172_ ),
    .Y(\soc/cpu/_04175_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08976_  (.A(\soc/cpu/decoded_imm_j[4] ),
    .B(\soc/cpu/_04162_ ),
    .Y(\soc/cpu/_04176_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_08977_  (.A1(\soc/cpu/_04150_ ),
    .A2(\soc/cpu/_04151_ ),
    .B1(\soc/cpu/_04162_ ),
    .B2(\soc/cpu/decoded_imm_j[4] ),
    .C1(\soc/cpu/_04152_ ),
    .Y(\soc/cpu/_04177_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08978_  (.A(\soc/cpu/_04176_ ),
    .B(\soc/cpu/_04177_ ),
    .Y(\soc/cpu/_04178_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08979_  (.A(\soc/cpu/_04175_ ),
    .B(\soc/cpu/_04178_ ),
    .Y(\soc/cpu/_04179_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_08980_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04172_ ),
    .B1(\soc/cpu/_04179_ ),
    .B2(\soc/cpu/_03312_ ),
    .Y(\soc/cpu/_04180_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08981_  (.A1(\soc/cpu/_04174_ ),
    .A2(\soc/cpu/_04180_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04181_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08982_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[5] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04172_ ),
    .C1(\soc/cpu/_04181_ ),
    .Y(\soc/cpu/_04182_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08983_  (.A(net132),
    .B(\soc/cpu/_04182_ ),
    .Y(\soc/cpu/_00348_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_08984_  (.A1(\soc/cpu/reg_next_pc[6] ),
    .A2(net161),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04183_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_08985_  (.A1(net161),
    .A2(\soc/cpu/_02159_ ),
    .B1(\soc/cpu/_04183_ ),
    .Y(\soc/cpu/_04184_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08986_  (.A(\soc/cpu/decoded_imm_j[5] ),
    .B(\soc/cpu/_04172_ ),
    .Y(\soc/cpu/_04185_ ));
 sky130_fd_sc_hd__o31a_1 \soc/cpu/_08987_  (.A1(\soc/cpu/_04176_ ),
    .A2(\soc/cpu/_04175_ ),
    .A3(\soc/cpu/_04177_ ),
    .B1(\soc/cpu/_04185_ ),
    .X(\soc/cpu/_04186_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08988_  (.A(\soc/cpu/decoded_imm_j[6] ),
    .B(\soc/cpu/_04184_ ),
    .Y(\soc/cpu/_04187_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_08989_  (.A1(\soc/cpu/_04186_ ),
    .A2(\soc/cpu/_04187_ ),
    .B1(\soc/cpu/_03312_ ),
    .Y(\soc/cpu/_04188_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_08990_  (.A1(\soc/cpu/_04186_ ),
    .A2(\soc/cpu/_04187_ ),
    .B1(\soc/cpu/_04188_ ),
    .X(\soc/cpu/_04189_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_08991_  (.A(\soc/cpu/_04156_ ),
    .B(\soc/cpu/_04162_ ),
    .C(\soc/cpu/_04172_ ),
    .D(\soc/cpu/_04184_ ),
    .Y(\soc/cpu/_04190_ ));
 sky130_fd_sc_hd__a31o_1 \soc/cpu/_08992_  (.A1(\soc/cpu/_04156_ ),
    .A2(\soc/cpu/_04162_ ),
    .A3(\soc/cpu/_04172_ ),
    .B1(\soc/cpu/_04184_ ),
    .X(\soc/cpu/_04191_ ));
 sky130_fd_sc_hd__a32oi_1 \soc/cpu/_08993_  (.A1(\soc/cpu/_04123_ ),
    .A2(\soc/cpu/_04190_ ),
    .A3(\soc/cpu/_04191_ ),
    .B1(\soc/cpu/_04131_ ),
    .B2(\soc/cpu/_04184_ ),
    .Y(\soc/cpu/_04192_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_08994_  (.A1(\soc/cpu/_04189_ ),
    .A2(\soc/cpu/_04192_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04193_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_08995_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[6] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04184_ ),
    .C1(\soc/cpu/_04193_ ),
    .Y(\soc/cpu/_04194_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_08996_  (.A(net131),
    .B(\soc/cpu/_04194_ ),
    .Y(\soc/cpu/_00349_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_08997_  (.A1(\soc/cpu/_02108_ ),
    .A2(net396),
    .B1(net161),
    .B2(\soc/cpu/_02164_ ),
    .C1(\soc/cpu/_01628_ ),
    .Y(\soc/cpu/_04195_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_08998_  (.A(\soc/cpu/_04190_ ),
    .B(\soc/cpu/_04195_ ),
    .Y(\soc/cpu/_04196_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_08999_  (.A(\soc/cpu/decoded_imm_j[6] ),
    .B(\soc/cpu/_04184_ ),
    .Y(\soc/cpu/_04197_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09000_  (.A1(\soc/cpu/_04186_ ),
    .A2(\soc/cpu/_04187_ ),
    .B1(\soc/cpu/_04197_ ),
    .X(\soc/cpu/_04198_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09001_  (.A(\soc/cpu/decoded_imm_j[7] ),
    .B(\soc/cpu/_04195_ ),
    .Y(\soc/cpu/_04199_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09002_  (.A(\soc/cpu/_04198_ ),
    .B(\soc/cpu/_04199_ ),
    .Y(\soc/cpu/_04200_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09003_  (.A(\soc/cpu/_04198_ ),
    .B(\soc/cpu/_04199_ ),
    .X(\soc/cpu/_04201_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09004_  (.A1(\soc/cpu/_04200_ ),
    .A2(\soc/cpu/_04201_ ),
    .B1(\soc/cpu/instr_jal ),
    .Y(\soc/cpu/_04202_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_09005_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04196_ ),
    .B1(\soc/cpu/_04202_ ),
    .C1(\soc/cpu/_00928_ ),
    .Y(\soc/cpu/_04203_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09007_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04195_ ),
    .B1(\soc/cpu/_04196_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04205_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09008_  (.A1(\soc/cpu/_04203_ ),
    .A2(\soc/cpu/_04205_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04206_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09009_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[7] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04195_ ),
    .C1(\soc/cpu/_04206_ ),
    .Y(\soc/cpu/_04207_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09010_  (.A(net131),
    .B(\soc/cpu/_04207_ ),
    .Y(\soc/cpu/_00350_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09011_  (.A1(\soc/cpu/reg_next_pc[8] ),
    .A2(net161),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04208_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09012_  (.A1(net161),
    .A2(\soc/cpu/_02170_ ),
    .B1(\soc/cpu/_04208_ ),
    .Y(\soc/cpu/_04209_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09013_  (.A_N(\soc/cpu/_04190_ ),
    .B(\soc/cpu/_04195_ ),
    .Y(\soc/cpu/_04210_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09014_  (.A(\soc/cpu/_04210_ ),
    .B(\soc/cpu/_04209_ ),
    .Y(\soc/cpu/_04211_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09015_  (.A(\soc/cpu/_03311_ ),
    .B(\soc/cpu/_04211_ ),
    .Y(\soc/cpu/_04212_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09016_  (.A1(\soc/cpu/decoded_imm_j[7] ),
    .A2(\soc/cpu/_04195_ ),
    .B1(\soc/cpu/_04200_ ),
    .Y(\soc/cpu/_04213_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09017_  (.A(\soc/cpu/decoded_imm_j[8] ),
    .B(\soc/cpu/_04209_ ),
    .Y(\soc/cpu/_04214_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09018_  (.A(\soc/cpu/decoded_imm_j[8] ),
    .B(\soc/cpu/_04209_ ),
    .Y(\soc/cpu/_04215_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09019_  (.A_N(\soc/cpu/_04214_ ),
    .B(\soc/cpu/_04215_ ),
    .Y(\soc/cpu/_04216_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09020_  (.A(\soc/cpu/_04213_ ),
    .B(\soc/cpu/_04216_ ),
    .Y(\soc/cpu/_04217_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09021_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04211_ ),
    .B1(\soc/cpu/_00928_ ),
    .Y(\soc/cpu/_04218_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09022_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04217_ ),
    .B1(\soc/cpu/_04218_ ),
    .Y(\soc/cpu/_04219_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09023_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04209_ ),
    .B1(\soc/cpu/_04219_ ),
    .Y(\soc/cpu/_04220_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09024_  (.A1(\soc/cpu/_04212_ ),
    .A2(\soc/cpu/_04220_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04221_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09025_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[8] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04209_ ),
    .C1(\soc/cpu/_04221_ ),
    .Y(\soc/cpu/_04222_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09026_  (.A(net131),
    .B(\soc/cpu/_04222_ ),
    .Y(\soc/cpu/_00351_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09029_  (.A1(net161),
    .A2(\soc/cpu/_02176_ ),
    .B1(net154),
    .Y(\soc/cpu/_04225_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/_09030_  (.A(\soc/cpu/_01639_ ),
    .B(\soc/cpu/_04225_ ),
    .Y(\soc/cpu/_04226_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09031_  (.A_N(\soc/cpu/_04210_ ),
    .B(\soc/cpu/_04209_ ),
    .Y(\soc/cpu/_04227_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09032_  (.A(\soc/cpu/_04227_ ),
    .B(\soc/cpu/_04226_ ),
    .Y(\soc/cpu/_04228_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09034_  (.A(\soc/cpu/decoded_imm_j[9] ),
    .B(\soc/cpu/_04226_ ),
    .Y(\soc/cpu/_04230_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09035_  (.A(\soc/cpu/decoded_imm_j[7] ),
    .B(\soc/cpu/_04195_ ),
    .Y(\soc/cpu/_04231_ ));
 sky130_fd_sc_hd__o211a_1 \soc/cpu/_09036_  (.A1(\soc/cpu/_04198_ ),
    .A2(\soc/cpu/_04199_ ),
    .B1(\soc/cpu/_04215_ ),
    .C1(\soc/cpu/_04231_ ),
    .X(\soc/cpu/_04232_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09037_  (.A(\soc/cpu/_04214_ ),
    .B(\soc/cpu/_04232_ ),
    .Y(\soc/cpu/_04233_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09038_  (.A(\soc/cpu/_04230_ ),
    .B(\soc/cpu/_04233_ ),
    .X(\soc/cpu/_04234_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09039_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04228_ ),
    .B1(\soc/cpu/_00928_ ),
    .Y(\soc/cpu/_04235_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09040_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04234_ ),
    .B1(\soc/cpu/_04235_ ),
    .Y(\soc/cpu/_04236_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09041_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04226_ ),
    .B1(\soc/cpu/_04228_ ),
    .B2(\soc/cpu/_03311_ ),
    .C1(\soc/cpu/_04236_ ),
    .Y(\soc/cpu/_04237_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09042_  (.A(\soc/cpu/_03994_ ),
    .B(\soc/cpu/_04237_ ),
    .Y(\soc/cpu/_04238_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09043_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[9] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04226_ ),
    .C1(\soc/cpu/_04238_ ),
    .Y(\soc/cpu/_04239_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09044_  (.A(net131),
    .B(\soc/cpu/_04239_ ),
    .Y(\soc/cpu/_00352_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09045_  (.A1(\soc/cpu/reg_next_pc[10] ),
    .A2(net161),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04240_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09046_  (.A1(net161),
    .A2(\soc/cpu/_02180_ ),
    .B1(\soc/cpu/_04240_ ),
    .Y(\soc/cpu/_04241_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09047_  (.A(\soc/cpu/decoded_imm_j[9] ),
    .B(\soc/cpu/_04226_ ),
    .Y(\soc/cpu/_04242_ ));
 sky130_fd_sc_hd__o31ai_2 \soc/cpu/_09048_  (.A1(\soc/cpu/_04214_ ),
    .A2(\soc/cpu/_04230_ ),
    .A3(\soc/cpu/_04232_ ),
    .B1(\soc/cpu/_04242_ ),
    .Y(\soc/cpu/_04243_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09049_  (.A(\soc/cpu/decoded_imm_j[10] ),
    .B(\soc/cpu/_04241_ ),
    .Y(\soc/cpu/_04244_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09050_  (.A(\soc/cpu/_04243_ ),
    .B(\soc/cpu/_04244_ ),
    .Y(\soc/cpu/_04245_ ));
 sky130_fd_sc_hd__and3b_1 \soc/cpu/_09051_  (.A_N(\soc/cpu/_04210_ ),
    .B(\soc/cpu/_04209_ ),
    .C(\soc/cpu/_04226_ ),
    .X(\soc/cpu/_04246_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09052_  (.A1(\soc/cpu/_04246_ ),
    .A2(\soc/cpu/_04241_ ),
    .B1(\soc/cpu/_04123_ ),
    .Y(\soc/cpu/_04247_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09053_  (.A1(\soc/cpu/_04246_ ),
    .A2(\soc/cpu/_04241_ ),
    .B1(\soc/cpu/_04247_ ),
    .Y(\soc/cpu/_04248_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_09054_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04241_ ),
    .B1(\soc/cpu/_04245_ ),
    .B2(\soc/cpu/_03312_ ),
    .C1(\soc/cpu/_04248_ ),
    .Y(\soc/cpu/_04249_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \soc/cpu/_09055_  (.A1_N(\soc/cpu/_00839_ ),
    .A2_N(\soc/cpu/reg_next_pc[10] ),
    .B1(\soc/cpu/_03994_ ),
    .B2(\soc/cpu/_04249_ ),
    .Y(\soc/cpu/_04250_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09056_  (.A1(\soc/cpu/_04114_ ),
    .A2(\soc/cpu/_04241_ ),
    .B1(\soc/cpu/_04250_ ),
    .Y(\soc/cpu/_04251_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09057_  (.A(net131),
    .B(\soc/cpu/_04251_ ),
    .Y(\soc/cpu/_00353_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09059_  (.A1(\soc/cpu/reg_next_pc[11] ),
    .A2(net161),
    .B1(net154),
    .Y(\soc/cpu/_04253_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_09060_  (.A1(\soc/cpu/_00709_ ),
    .A2(\soc/cpu/_02185_ ),
    .B1(\soc/cpu/_04253_ ),
    .Y(\soc/cpu/_04254_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09061_  (.A(\soc/cpu/_04246_ ),
    .B(\soc/cpu/_04241_ ),
    .Y(\soc/cpu/_04255_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09062_  (.A(\soc/cpu/_04255_ ),
    .B(\soc/cpu/_04254_ ),
    .Y(\soc/cpu/_04256_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09063_  (.A(\soc/cpu/decoded_imm_j[11] ),
    .B(\soc/cpu/_04254_ ),
    .Y(\soc/cpu/_04257_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09064_  (.A(\soc/cpu/_04257_ ),
    .Y(\soc/cpu/_04258_ ));
 sky130_fd_sc_hd__maj3_2 \soc/cpu/_09065_  (.A(\soc/cpu/decoded_imm_j[10] ),
    .B(\soc/cpu/_04243_ ),
    .C(\soc/cpu/_04241_ ),
    .X(\soc/cpu/_04259_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09066_  (.A(\soc/cpu/_04258_ ),
    .B(\soc/cpu/_04259_ ),
    .Y(\soc/cpu/_04260_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09067_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04260_ ),
    .B1(\soc/cpu/_03993_ ),
    .Y(\soc/cpu/_04261_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09068_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04256_ ),
    .B1(\soc/cpu/_04261_ ),
    .Y(\soc/cpu/_04262_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09069_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04254_ ),
    .B1(\soc/cpu/_04256_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04263_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09070_  (.A1(\soc/cpu/_04262_ ),
    .A2(\soc/cpu/_04263_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04264_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09071_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[11] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04254_ ),
    .C1(\soc/cpu/_04264_ ),
    .Y(\soc/cpu/_04265_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09072_  (.A(net131),
    .B(\soc/cpu/_04265_ ),
    .Y(\soc/cpu/_00354_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09073_  (.A1(\soc/cpu/reg_next_pc[12] ),
    .A2(net161),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04266_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09074_  (.A1(net161),
    .A2(\soc/cpu/_02190_ ),
    .B1(\soc/cpu/_04266_ ),
    .Y(\soc/cpu/_04267_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09075_  (.A(\soc/cpu/_03300_ ),
    .B(\soc/cpu/_04267_ ),
    .Y(\soc/cpu/_04268_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09076_  (.A(\soc/cpu/_04246_ ),
    .B(\soc/cpu/_04241_ ),
    .C(\soc/cpu/_04254_ ),
    .Y(\soc/cpu/_04269_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09077_  (.A(\soc/cpu/_04269_ ),
    .B(\soc/cpu/_04267_ ),
    .Y(\soc/cpu/_04270_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09078_  (.A(\soc/cpu/decoded_imm_j[11] ),
    .B(\soc/cpu/_04254_ ),
    .X(\soc/cpu/_04271_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_09079_  (.A1(\soc/cpu/_04258_ ),
    .A2(\soc/cpu/_04259_ ),
    .B1(\soc/cpu/_04271_ ),
    .X(\soc/cpu/_04272_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09080_  (.A(\soc/cpu/decoded_imm_j[12] ),
    .B(\soc/cpu/_04267_ ),
    .Y(\soc/cpu/_04273_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09081_  (.A(\soc/cpu/decoded_imm_j[12] ),
    .B(\soc/cpu/_04267_ ),
    .Y(\soc/cpu/_04274_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09082_  (.A(\soc/cpu/_04274_ ),
    .Y(\soc/cpu/_04275_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09083_  (.A(\soc/cpu/_04273_ ),
    .B(\soc/cpu/_04275_ ),
    .Y(\soc/cpu/_04276_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09084_  (.A(\soc/cpu/_04272_ ),
    .B(\soc/cpu/_04276_ ),
    .Y(\soc/cpu/_04277_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09085_  (.A(\soc/cpu/_00926_ ),
    .B(\soc/cpu/_04277_ ),
    .Y(\soc/cpu/_04278_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09086_  (.A1(\soc/cpu/_00746_ ),
    .A2(\soc/cpu/_04267_ ),
    .B1(\soc/cpu/_04270_ ),
    .B2(\soc/cpu/_00818_ ),
    .C1(\soc/cpu/_04278_ ),
    .Y(\soc/cpu/_04279_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \soc/cpu/_09087_  (.A1_N(\soc/cpu/_00924_ ),
    .A2_N(\soc/cpu/_04279_ ),
    .B1(\soc/cpu/_04270_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04280_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09088_  (.A1(\soc/cpu/_04268_ ),
    .A2(\soc/cpu/_04280_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04281_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09089_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[12] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04267_ ),
    .C1(\soc/cpu/_04281_ ),
    .Y(\soc/cpu/_04282_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09090_  (.A(net131),
    .B(\soc/cpu/_04282_ ),
    .Y(\soc/cpu/_00355_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09091_  (.A(\soc/cpu/_01659_ ),
    .B(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04283_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09092_  (.A1(net161),
    .A2(\soc/cpu/_02193_ ),
    .B1(\soc/cpu/_04283_ ),
    .Y(\soc/cpu/_04284_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09093_  (.A(\soc/cpu/_04246_ ),
    .B(\soc/cpu/_04241_ ),
    .C(\soc/cpu/_04254_ ),
    .D(\soc/cpu/_04267_ ),
    .Y(\soc/cpu/_04285_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09094_  (.A(\soc/cpu/_04285_ ),
    .B(\soc/cpu/_04284_ ),
    .Y(\soc/cpu/_04286_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_09095_  (.A(\soc/cpu/decoded_imm_j[13] ),
    .B(\soc/cpu/_04284_ ),
    .Y(\soc/cpu/_04287_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_09096_  (.A1(\soc/cpu/_04258_ ),
    .A2(\soc/cpu/_04259_ ),
    .B1(\soc/cpu/_04275_ ),
    .C1(\soc/cpu/_04271_ ),
    .Y(\soc/cpu/_04288_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09097_  (.A(\soc/cpu/_04273_ ),
    .B(\soc/cpu/_04288_ ),
    .Y(\soc/cpu/_04289_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09098_  (.A(\soc/cpu/_04287_ ),
    .B(\soc/cpu/_04289_ ),
    .X(\soc/cpu/_04290_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09099_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04290_ ),
    .B1(\soc/cpu/_03993_ ),
    .Y(\soc/cpu/_04291_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09100_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04286_ ),
    .B1(\soc/cpu/_04291_ ),
    .Y(\soc/cpu/_04292_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09101_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04284_ ),
    .B1(\soc/cpu/_04286_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04293_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09103_  (.A1(\soc/cpu/_04292_ ),
    .A2(\soc/cpu/_04293_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04295_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09104_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[13] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04284_ ),
    .C1(\soc/cpu/_04295_ ),
    .Y(\soc/cpu/_04296_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09105_  (.A(net131),
    .B(\soc/cpu/_04296_ ),
    .Y(\soc/cpu/_00356_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09106_  (.A(\soc/cpu/_00709_ ),
    .B(\soc/cpu/_02199_ ),
    .Y(\soc/cpu/_04297_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09107_  (.A1(\soc/cpu/reg_next_pc[14] ),
    .A2(net161),
    .B1(net154),
    .B2(\soc/cpu/_04297_ ),
    .X(\soc/cpu/_04298_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09108_  (.A(\soc/cpu/decoded_imm_j[13] ),
    .B(\soc/cpu/_04284_ ),
    .Y(\soc/cpu/_04299_ ));
 sky130_fd_sc_hd__o31a_1 \soc/cpu/_09109_  (.A1(\soc/cpu/_04273_ ),
    .A2(\soc/cpu/_04287_ ),
    .A3(\soc/cpu/_04288_ ),
    .B1(\soc/cpu/_04299_ ),
    .X(\soc/cpu/_04300_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09110_  (.A(\soc/cpu/decoded_imm_j[14] ),
    .B(\soc/cpu/_04298_ ),
    .Y(\soc/cpu/_04301_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_09111_  (.A(\soc/cpu/decoded_imm_j[14] ),
    .B(\soc/cpu/_04298_ ),
    .X(\soc/cpu/_04302_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09112_  (.A(\soc/cpu/_04301_ ),
    .B(\soc/cpu/_04302_ ),
    .Y(\soc/cpu/_04303_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09113_  (.A(\soc/cpu/_04300_ ),
    .B(\soc/cpu/_04303_ ),
    .Y(\soc/cpu/_04304_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09114_  (.A(\soc/cpu/_00926_ ),
    .B(\soc/cpu/_04304_ ),
    .Y(\soc/cpu/_04305_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/_09115_  (.A1(\soc/cpu/reg_next_pc[14] ),
    .A2(net161),
    .B1(net154),
    .B2(\soc/cpu/_04297_ ),
    .Y(\soc/cpu/_04306_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09116_  (.A_N(\soc/cpu/_04285_ ),
    .B(\soc/cpu/_04284_ ),
    .Y(\soc/cpu/_04307_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09117_  (.A(\soc/cpu/_04307_ ),
    .B(\soc/cpu/_04306_ ),
    .Y(\soc/cpu/_04308_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_09118_  (.A1(\soc/cpu/decoder_trigger ),
    .A2(\soc/cpu/_04306_ ),
    .B1(\soc/cpu/_04308_ ),
    .B2(\soc/cpu/_03322_ ),
    .Y(\soc/cpu/_04309_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09119_  (.A1(\soc/cpu/_04305_ ),
    .A2(\soc/cpu/_04309_ ),
    .B1(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04310_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09120_  (.A(\soc/cpu/_03403_ ),
    .B(\soc/cpu/_04308_ ),
    .Y(\soc/cpu/_04311_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09121_  (.A1(\soc/cpu/_03300_ ),
    .A2(\soc/cpu/_04298_ ),
    .B1(\soc/cpu/_04311_ ),
    .Y(\soc/cpu/_04312_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09122_  (.A1(\soc/cpu/_04310_ ),
    .A2(\soc/cpu/_04312_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04313_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09123_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[14] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04298_ ),
    .C1(\soc/cpu/_04313_ ),
    .Y(\soc/cpu/_04314_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09124_  (.A(net131),
    .B(\soc/cpu/_04314_ ),
    .Y(\soc/cpu/_00357_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09125_  (.A1(\soc/cpu/reg_next_pc[15] ),
    .A2(net161),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04315_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09126_  (.A1(net161),
    .A2(\soc/cpu/_02204_ ),
    .B1(\soc/cpu/_04315_ ),
    .Y(\soc/cpu/_04316_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09127_  (.A_N(\soc/cpu/_04300_ ),
    .B(\soc/cpu/_04302_ ),
    .Y(\soc/cpu/_04317_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_09128_  (.A(\soc/cpu/decoded_imm_j[15] ),
    .B(\soc/cpu/_04316_ ),
    .X(\soc/cpu/_04318_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09129_  (.A(\soc/cpu/decoded_imm_j[15] ),
    .B(\soc/cpu/_04316_ ),
    .Y(\soc/cpu/_04319_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09130_  (.A(\soc/cpu/_04318_ ),
    .B(\soc/cpu/_04319_ ),
    .Y(\soc/cpu/_04320_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09131_  (.A1(\soc/cpu/_04301_ ),
    .A2(\soc/cpu/_04317_ ),
    .B1(\soc/cpu/_04320_ ),
    .Y(\soc/cpu/_04321_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09132_  (.A(\soc/cpu/_04301_ ),
    .B(\soc/cpu/_04317_ ),
    .C(\soc/cpu/_04320_ ),
    .Y(\soc/cpu/_04322_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_09133_  (.A_N(\soc/cpu/_04321_ ),
    .B(\soc/cpu/_04322_ ),
    .C(\soc/cpu/_03312_ ),
    .Y(\soc/cpu/_04323_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09134_  (.A(\soc/cpu/_04307_ ),
    .B(\soc/cpu/_04306_ ),
    .Y(\soc/cpu/_04324_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09135_  (.A(\soc/cpu/_04324_ ),
    .B(\soc/cpu/_04316_ ),
    .X(\soc/cpu/_04325_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09136_  (.A(\soc/cpu/_03311_ ),
    .B(\soc/cpu/_04325_ ),
    .Y(\soc/cpu/_04326_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09137_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04316_ ),
    .B1(\soc/cpu/_04325_ ),
    .B2(\soc/cpu/_03323_ ),
    .Y(\soc/cpu/_04327_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/cpu/_09138_  (.A1(\soc/cpu/_04323_ ),
    .A2(\soc/cpu/_04326_ ),
    .A3(\soc/cpu/_04327_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04328_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09139_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[15] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04316_ ),
    .C1(\soc/cpu/_04328_ ),
    .Y(\soc/cpu/_04329_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09140_  (.A(net131),
    .B(\soc/cpu/_04329_ ),
    .Y(\soc/cpu/_00358_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09142_  (.A1(\soc/cpu/reg_next_pc[16] ),
    .A2(net161),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04331_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09143_  (.A1(net161),
    .A2(\soc/cpu/_02207_ ),
    .B1(\soc/cpu/_04331_ ),
    .Y(\soc/cpu/_04332_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09144_  (.A(\soc/cpu/_04114_ ),
    .B(\soc/cpu/_04332_ ),
    .Y(\soc/cpu/_04333_ ));
 sky130_fd_sc_hd__nor3b_2 \soc/cpu/_09145_  (.A(\soc/cpu/_04307_ ),
    .B(\soc/cpu/_04306_ ),
    .C_N(\soc/cpu/_04316_ ),
    .Y(\soc/cpu/_04334_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09146_  (.A(\soc/cpu/_04334_ ),
    .B(\soc/cpu/_04332_ ),
    .X(\soc/cpu/_04335_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09147_  (.A(\soc/cpu/decoded_imm_j[15] ),
    .B(\soc/cpu/_04316_ ),
    .X(\soc/cpu/_04336_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09148_  (.A(\soc/cpu/decoded_imm_j[16] ),
    .B(\soc/cpu/_04332_ ),
    .Y(\soc/cpu/_04337_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09149_  (.A(\soc/cpu/_04337_ ),
    .Y(\soc/cpu/_04338_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09150_  (.A(\soc/cpu/_04336_ ),
    .B(\soc/cpu/_04321_ ),
    .C(\soc/cpu/_04338_ ),
    .Y(\soc/cpu/_04339_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09151_  (.A1(\soc/cpu/decoded_imm_j[16] ),
    .A2(\soc/cpu/_04332_ ),
    .B1(\soc/cpu/_04339_ ),
    .Y(\soc/cpu/_04340_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09152_  (.A(\soc/cpu/decoded_imm_j[16] ),
    .B(\soc/cpu/_04332_ ),
    .Y(\soc/cpu/_04341_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_09153_  (.A1(\soc/cpu/_04336_ ),
    .A2(\soc/cpu/_04321_ ),
    .B1(\soc/cpu/_04341_ ),
    .B2(\soc/cpu/_04338_ ),
    .Y(\soc/cpu/_04342_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09154_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04335_ ),
    .B1(\soc/cpu/_00928_ ),
    .Y(\soc/cpu/_04343_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09155_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04340_ ),
    .A3(\soc/cpu/_04342_ ),
    .B1(\soc/cpu/_04343_ ),
    .Y(\soc/cpu/_04344_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/_09156_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04332_ ),
    .B1(\soc/cpu/_04335_ ),
    .B2(\soc/cpu/_03311_ ),
    .C1(\soc/cpu/_04344_ ),
    .Y(\soc/cpu/_04345_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09157_  (.A(\soc/cpu/_03994_ ),
    .B(\soc/cpu/_04345_ ),
    .Y(\soc/cpu/_04346_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09158_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[16] ),
    .B1(\soc/cpu/_04346_ ),
    .Y(\soc/cpu/_04347_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09159_  (.A1(\soc/cpu/_04333_ ),
    .A2(\soc/cpu/_04347_ ),
    .B1(net131),
    .Y(\soc/cpu/_00359_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09160_  (.A1(\soc/cpu/reg_next_pc[17] ),
    .A2(net161),
    .B1(net154),
    .Y(\soc/cpu/_04348_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_09161_  (.A1(\soc/cpu/_00709_ ),
    .A2(\soc/cpu/_02213_ ),
    .B1(\soc/cpu/_04348_ ),
    .Y(\soc/cpu/_04349_ ));
 sky130_fd_sc_hd__o311ai_2 \soc/cpu/_09162_  (.A1(\soc/cpu/_04273_ ),
    .A2(\soc/cpu/_04287_ ),
    .A3(\soc/cpu/_04288_ ),
    .B1(\soc/cpu/_04301_ ),
    .C1(\soc/cpu/_04299_ ),
    .Y(\soc/cpu/_04350_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09163_  (.A1(\soc/cpu/_04302_ ),
    .A2(\soc/cpu/_04318_ ),
    .A3(\soc/cpu/_04350_ ),
    .B1(\soc/cpu/_04336_ ),
    .Y(\soc/cpu/_04351_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09164_  (.A(\soc/cpu/decoded_imm_j[17] ),
    .B(\soc/cpu/_04349_ ),
    .Y(\soc/cpu/_04352_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/cpu/_09165_  (.A1(\soc/cpu/_04351_ ),
    .A2(\soc/cpu/_04337_ ),
    .B1(\soc/cpu/_04352_ ),
    .C1(\soc/cpu/_04341_ ),
    .Y(\soc/cpu/_04353_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09166_  (.A1(\soc/cpu/_04341_ ),
    .A2(\soc/cpu/_04339_ ),
    .B1(\soc/cpu/_04352_ ),
    .Y(\soc/cpu/_04354_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/cpu/_09167_  (.A_N(\soc/cpu/_04353_ ),
    .B(\soc/cpu/_04354_ ),
    .C(\soc/cpu/_03312_ ),
    .Y(\soc/cpu/_04355_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_09168_  (.A1(\soc/cpu/_04334_ ),
    .A2(\soc/cpu/_04332_ ),
    .B1(\soc/cpu/_04349_ ),
    .X(\soc/cpu/_04356_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09169_  (.A(\soc/cpu/_04334_ ),
    .B(\soc/cpu/_04332_ ),
    .C(\soc/cpu/_04349_ ),
    .Y(\soc/cpu/_04357_ ));
 sky130_fd_sc_hd__a32oi_1 \soc/cpu/_09170_  (.A1(\soc/cpu/_04123_ ),
    .A2(\soc/cpu/_04356_ ),
    .A3(\soc/cpu/_04357_ ),
    .B1(\soc/cpu/_04131_ ),
    .B2(\soc/cpu/_04349_ ),
    .Y(\soc/cpu/_04358_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09171_  (.A1(\soc/cpu/_04355_ ),
    .A2(\soc/cpu/_04358_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04359_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09172_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[17] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04349_ ),
    .C1(\soc/cpu/_04359_ ),
    .Y(\soc/cpu/_04360_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09173_  (.A(net131),
    .B(\soc/cpu/_04360_ ),
    .Y(\soc/cpu/_00360_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09174_  (.A1(\soc/cpu/reg_next_pc[18] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04361_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09175_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02218_ ),
    .B1(\soc/cpu/_04361_ ),
    .Y(\soc/cpu/_04362_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09176_  (.A1(\soc/cpu/decoded_imm_j[17] ),
    .A2(\soc/cpu/_04349_ ),
    .B1(\soc/cpu/_04353_ ),
    .Y(\soc/cpu/_04363_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09177_  (.A(\soc/cpu/decoded_imm_j[18] ),
    .B(\soc/cpu/_04362_ ),
    .Y(\soc/cpu/_04364_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09178_  (.A(\soc/cpu/_04363_ ),
    .B(\soc/cpu/_04364_ ),
    .Y(\soc/cpu/_04365_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09179_  (.A(\soc/cpu/_00926_ ),
    .B(\soc/cpu/_04365_ ),
    .Y(\soc/cpu/_04366_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09180_  (.A(\soc/cpu/_04362_ ),
    .Y(\soc/cpu/_04367_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_09181_  (.A(\soc/cpu/_04334_ ),
    .B(\soc/cpu/_04332_ ),
    .C(\soc/cpu/_04349_ ),
    .D(\soc/cpu/_04362_ ),
    .Y(\soc/cpu/_04368_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09182_  (.A(\soc/cpu/_04357_ ),
    .B(\soc/cpu/_04367_ ),
    .Y(\soc/cpu/_04369_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09183_  (.A(\soc/cpu/_04368_ ),
    .B(\soc/cpu/_04369_ ),
    .Y(\soc/cpu/_04370_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_09184_  (.A1(\soc/cpu/decoder_trigger ),
    .A2(\soc/cpu/_04367_ ),
    .B1(\soc/cpu/_04370_ ),
    .B2(\soc/cpu/_03322_ ),
    .Y(\soc/cpu/_04371_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09185_  (.A1(\soc/cpu/_04366_ ),
    .A2(\soc/cpu/_04371_ ),
    .B1(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04372_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09186_  (.A(\soc/cpu/_03403_ ),
    .B(\soc/cpu/_04370_ ),
    .Y(\soc/cpu/_04373_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09187_  (.A1(\soc/cpu/_03300_ ),
    .A2(\soc/cpu/_04362_ ),
    .B1(\soc/cpu/_04373_ ),
    .Y(\soc/cpu/_04374_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09188_  (.A1(\soc/cpu/_04372_ ),
    .A2(\soc/cpu/_04374_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04375_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09189_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[18] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04362_ ),
    .C1(\soc/cpu/_04375_ ),
    .Y(\soc/cpu/_04376_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09190_  (.A(net131),
    .B(\soc/cpu/_04376_ ),
    .Y(\soc/cpu/_00361_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \soc/cpu/_09191_  (.A1_N(\soc/cpu/_01683_ ),
    .A2_N(net154),
    .B1(\soc/cpu/_02223_ ),
    .B2(\soc/cpu/_00709_ ),
    .Y(\soc/cpu/_04377_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09192_  (.A(\soc/cpu/_04368_ ),
    .B(\soc/cpu/_04377_ ),
    .Y(\soc/cpu/_04378_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_09193_  (.A(\soc/cpu/decoded_imm_j[19] ),
    .B(\soc/cpu/_04377_ ),
    .Y(\soc/cpu/_04379_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09194_  (.A(\soc/cpu/decoded_imm_j[18] ),
    .B(\soc/cpu/_04362_ ),
    .Y(\soc/cpu/_04380_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/cpu/_09195_  (.A1(\soc/cpu/decoded_imm_j[17] ),
    .A2(\soc/cpu/_04349_ ),
    .B1(\soc/cpu/_04362_ ),
    .B2(\soc/cpu/decoded_imm_j[18] ),
    .C1(\soc/cpu/_04353_ ),
    .Y(\soc/cpu/_04381_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09196_  (.A(\soc/cpu/_04380_ ),
    .B(\soc/cpu/_04381_ ),
    .Y(\soc/cpu/_04382_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09197_  (.A(\soc/cpu/_04379_ ),
    .B(\soc/cpu/_04382_ ),
    .X(\soc/cpu/_04383_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09198_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04383_ ),
    .B1(\soc/cpu/_03993_ ),
    .Y(\soc/cpu/_04384_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09199_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04378_ ),
    .B1(\soc/cpu/_04384_ ),
    .Y(\soc/cpu/_04385_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09200_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04377_ ),
    .B1(\soc/cpu/_04378_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04386_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09201_  (.A1(\soc/cpu/_04385_ ),
    .A2(\soc/cpu/_04386_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04387_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09202_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[19] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04377_ ),
    .C1(\soc/cpu/_04387_ ),
    .Y(\soc/cpu/_04388_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09203_  (.A(net131),
    .B(\soc/cpu/_04388_ ),
    .Y(\soc/cpu/_00362_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09204_  (.A1(\soc/cpu/reg_next_pc[20] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04389_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09205_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02228_ ),
    .B1(\soc/cpu/_04389_ ),
    .Y(\soc/cpu/_04390_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09206_  (.A_N(\soc/cpu/_04368_ ),
    .B(\soc/cpu/_04377_ ),
    .Y(\soc/cpu/_04391_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09207_  (.A(\soc/cpu/_04391_ ),
    .B(\soc/cpu/_04390_ ),
    .Y(\soc/cpu/_04392_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09208_  (.A(\soc/cpu/decoded_imm_j[19] ),
    .B(\soc/cpu/_04377_ ),
    .Y(\soc/cpu/_04393_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_09209_  (.A1(\soc/cpu/_04380_ ),
    .A2(\soc/cpu/_04379_ ),
    .A3(\soc/cpu/_04381_ ),
    .B1(\soc/cpu/_04393_ ),
    .Y(\soc/cpu/_04394_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09210_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04390_ ),
    .Y(\soc/cpu/_04395_ ));
 sky130_fd_sc_hd__or2_0 \soc/cpu/_09211_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04390_ ),
    .X(\soc/cpu/_04396_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09212_  (.A(\soc/cpu/_04395_ ),
    .B(\soc/cpu/_04396_ ),
    .Y(\soc/cpu/_04397_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09213_  (.A(\soc/cpu/_04394_ ),
    .B(\soc/cpu/_04397_ ),
    .X(\soc/cpu/_04398_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09214_  (.A(\soc/cpu/_00926_ ),
    .B(\soc/cpu/_04398_ ),
    .Y(\soc/cpu/_04399_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09215_  (.A1(\soc/cpu/_00746_ ),
    .A2(\soc/cpu/_04390_ ),
    .B1(\soc/cpu/_04392_ ),
    .B2(\soc/cpu/_00818_ ),
    .C1(\soc/cpu/_04399_ ),
    .Y(\soc/cpu/_04400_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09216_  (.A(\soc/cpu/_00924_ ),
    .B(\soc/cpu/_04400_ ),
    .Y(\soc/cpu/_04401_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09217_  (.A1(\soc/cpu/_03300_ ),
    .A2(\soc/cpu/_04390_ ),
    .B1(\soc/cpu/_04392_ ),
    .B2(\soc/cpu/_03311_ ),
    .C1(\soc/cpu/_04401_ ),
    .Y(\soc/cpu/_04402_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09218_  (.A(\soc/cpu/_04114_ ),
    .B(\soc/cpu/_04390_ ),
    .Y(\soc/cpu/_04403_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09219_  (.A(\soc/cpu/_00839_ ),
    .B(\soc/cpu/reg_next_pc[20] ),
    .Y(\soc/cpu/_04404_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/cpu/_09220_  (.A1(\soc/cpu/_03994_ ),
    .A2(\soc/cpu/_04402_ ),
    .B1(\soc/cpu/_04403_ ),
    .C1(\soc/cpu/_04404_ ),
    .D1(_074_),
    .Y(\soc/cpu/_00363_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09222_  (.A(\soc/cpu/_01693_ ),
    .B(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04406_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09223_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02231_ ),
    .B1(\soc/cpu/_04406_ ),
    .Y(\soc/cpu/_04407_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_09224_  (.A(\soc/cpu/_04391_ ),
    .B_N(\soc/cpu/_04390_ ),
    .Y(\soc/cpu/_04408_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09225_  (.A(\soc/cpu/_04408_ ),
    .B(\soc/cpu/_04407_ ),
    .X(\soc/cpu/_04409_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09226_  (.A(\soc/cpu/_02484_ ),
    .B(\soc/cpu/_04407_ ),
    .Y(\soc/cpu/_04410_ ));
 sky130_fd_sc_hd__o311ai_2 \soc/cpu/_09227_  (.A1(\soc/cpu/_04380_ ),
    .A2(\soc/cpu/_04379_ ),
    .A3(\soc/cpu/_04381_ ),
    .B1(\soc/cpu/_04395_ ),
    .C1(\soc/cpu/_04393_ ),
    .Y(\soc/cpu/_04411_ ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_09228_  (.A(\soc/cpu/_04396_ ),
    .B(\soc/cpu/_04410_ ),
    .C(\soc/cpu/_04411_ ),
    .X(\soc/cpu/_04412_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09229_  (.A1(\soc/cpu/_04396_ ),
    .A2(\soc/cpu/_04411_ ),
    .B1(\soc/cpu/_04410_ ),
    .Y(\soc/cpu/_04413_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09230_  (.A1(\soc/cpu/_04412_ ),
    .A2(\soc/cpu/_04413_ ),
    .B1(\soc/cpu/instr_jal ),
    .Y(\soc/cpu/_04414_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/cpu/_09231_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04409_ ),
    .B1(\soc/cpu/_04414_ ),
    .C1(\soc/cpu/_00928_ ),
    .Y(\soc/cpu/_04415_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09232_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04407_ ),
    .B1(\soc/cpu/_04409_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04416_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09233_  (.A1(\soc/cpu/_04415_ ),
    .A2(\soc/cpu/_04416_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04417_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09234_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[21] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04407_ ),
    .C1(\soc/cpu/_04417_ ),
    .Y(\soc/cpu/_04418_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09235_  (.A(net131),
    .B(\soc/cpu/_04418_ ),
    .Y(\soc/cpu/_00364_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09236_  (.A(\soc/cpu/_01699_ ),
    .B(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04419_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09237_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02237_ ),
    .B1(\soc/cpu/_04419_ ),
    .Y(\soc/cpu/_04420_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09239_  (.A(\soc/cpu/_04420_ ),
    .SLEEP(\soc/cpu/decoder_trigger ),
    .X(\soc/cpu/_04422_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09240_  (.A1(\soc/cpu/decoded_imm_j[20] ),
    .A2(\soc/cpu/_04407_ ),
    .B1(\soc/cpu/_04412_ ),
    .Y(\soc/cpu/_04423_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/cpu/_09241_  (.A(\soc/cpu/_02484_ ),
    .B(\soc/cpu/_04420_ ),
    .Y(\soc/cpu/_04424_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09242_  (.A(\soc/cpu/_04423_ ),
    .B(\soc/cpu/_04424_ ),
    .X(\soc/cpu/_04425_ ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_09243_  (.A(\soc/cpu/_04408_ ),
    .B(\soc/cpu/_04407_ ),
    .X(\soc/cpu/_04426_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09244_  (.A(\soc/cpu/_04426_ ),
    .B(\soc/cpu/_04420_ ),
    .Y(\soc/cpu/_04427_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_09245_  (.A1(\soc/cpu/_00926_ ),
    .A2(\soc/cpu/_04425_ ),
    .B1(\soc/cpu/_04427_ ),
    .B2(\soc/cpu/_03322_ ),
    .Y(\soc/cpu/_04428_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09246_  (.A1(\soc/cpu/_04422_ ),
    .A2(\soc/cpu/_04428_ ),
    .B1(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04429_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09247_  (.A(\soc/cpu/_03403_ ),
    .B(\soc/cpu/_04427_ ),
    .Y(\soc/cpu/_04430_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09248_  (.A1(\soc/cpu/_03300_ ),
    .A2(\soc/cpu/_04420_ ),
    .B1(\soc/cpu/_04430_ ),
    .Y(\soc/cpu/_04431_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09249_  (.A1(\soc/cpu/_04429_ ),
    .A2(\soc/cpu/_04431_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04432_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09250_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[22] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04420_ ),
    .C1(\soc/cpu/_04432_ ),
    .Y(\soc/cpu/_04433_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09251_  (.A(net131),
    .B(\soc/cpu/_04433_ ),
    .Y(\soc/cpu/_00365_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09252_  (.A1(\soc/cpu/reg_next_pc[23] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04434_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09253_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02242_ ),
    .B1(\soc/cpu/_04434_ ),
    .Y(\soc/cpu/_04435_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09254_  (.A(\soc/cpu/_04114_ ),
    .B(\soc/cpu/_04435_ ),
    .Y(\soc/cpu/_04436_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09255_  (.A(\soc/cpu/_04426_ ),
    .B(\soc/cpu/_04420_ ),
    .Y(\soc/cpu/_04437_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09256_  (.A(\soc/cpu/_04437_ ),
    .B(\soc/cpu/_04435_ ),
    .Y(\soc/cpu/_04438_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09257_  (.A(\soc/cpu/_03311_ ),
    .B(\soc/cpu/_04438_ ),
    .Y(\soc/cpu/_04439_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09258_  (.A(\soc/cpu/_04131_ ),
    .B(\soc/cpu/_04435_ ),
    .Y(\soc/cpu/_04440_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09259_  (.A1(\soc/cpu/_04407_ ),
    .A2(\soc/cpu/_04420_ ),
    .B1(\soc/cpu/decoded_imm_j[20] ),
    .Y(\soc/cpu/_04441_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09260_  (.A(\soc/cpu/_04412_ ),
    .B(\soc/cpu/_04424_ ),
    .Y(\soc/cpu/_04442_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09261_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04435_ ),
    .Y(\soc/cpu/_04443_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09262_  (.A1(\soc/cpu/_04441_ ),
    .A2(\soc/cpu/_04442_ ),
    .B1(\soc/cpu/_04443_ ),
    .Y(\soc/cpu/_04444_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09263_  (.A(\soc/cpu/_04441_ ),
    .B(\soc/cpu/_04442_ ),
    .C(\soc/cpu/_04443_ ),
    .Y(\soc/cpu/_04445_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09264_  (.A_N(\soc/cpu/_04444_ ),
    .B(\soc/cpu/_04445_ ),
    .Y(\soc/cpu/_04446_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09265_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04446_ ),
    .B1(\soc/cpu/_03993_ ),
    .Y(\soc/cpu/_04447_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09266_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04438_ ),
    .B1(\soc/cpu/_04447_ ),
    .Y(\soc/cpu/_04448_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09267_  (.A1(\soc/cpu/_04439_ ),
    .A2(\soc/cpu/_04440_ ),
    .A3(\soc/cpu/_04448_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04449_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09268_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[23] ),
    .B1(\soc/cpu/_04449_ ),
    .Y(\soc/cpu/_04450_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09269_  (.A1(\soc/cpu/_04436_ ),
    .A2(\soc/cpu/_04450_ ),
    .B1(net131),
    .Y(\soc/cpu/_00366_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09270_  (.A1(\soc/cpu/reg_next_pc[24] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04451_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09271_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02245_ ),
    .B1(\soc/cpu/_04451_ ),
    .Y(\soc/cpu/_04452_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09272_  (.A(\soc/cpu/_04452_ ),
    .SLEEP(\soc/cpu/decoder_trigger ),
    .X(\soc/cpu/_04453_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09273_  (.A1(\soc/cpu/decoded_imm_j[20] ),
    .A2(\soc/cpu/_04435_ ),
    .B1(\soc/cpu/_04444_ ),
    .Y(\soc/cpu/_04454_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09274_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04452_ ),
    .Y(\soc/cpu/_04455_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09275_  (.A(\soc/cpu/_04454_ ),
    .B(\soc/cpu/_04455_ ),
    .Y(\soc/cpu/_04456_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_09276_  (.A(\soc/cpu/_04426_ ),
    .B(\soc/cpu/_04420_ ),
    .C(\soc/cpu/_04435_ ),
    .D(\soc/cpu/_04452_ ),
    .Y(\soc/cpu/_04457_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09277_  (.A1(\soc/cpu/_04426_ ),
    .A2(\soc/cpu/_04420_ ),
    .A3(\soc/cpu/_04435_ ),
    .B1(\soc/cpu/_04452_ ),
    .Y(\soc/cpu/_04458_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09278_  (.A(\soc/cpu/_04457_ ),
    .SLEEP(\soc/cpu/_04458_ ),
    .X(\soc/cpu/_04459_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09279_  (.A(\soc/cpu/_00818_ ),
    .B(\soc/cpu/_04459_ ),
    .Y(\soc/cpu/_04460_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09280_  (.A1(\soc/cpu/_00926_ ),
    .A2(\soc/cpu/_04456_ ),
    .B1(\soc/cpu/_04460_ ),
    .Y(\soc/cpu/_04461_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09281_  (.A1(\soc/cpu/_04453_ ),
    .A2(\soc/cpu/_04461_ ),
    .B1(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04462_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09282_  (.A1(\soc/cpu/_03300_ ),
    .A2(\soc/cpu/_04452_ ),
    .B1(\soc/cpu/_04459_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04463_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09283_  (.A1(\soc/cpu/_04462_ ),
    .A2(\soc/cpu/_04463_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04464_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09284_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[24] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04452_ ),
    .C1(\soc/cpu/_04464_ ),
    .Y(\soc/cpu/_04465_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09285_  (.A(net131),
    .B(\soc/cpu/_04465_ ),
    .Y(\soc/cpu/_00367_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09286_  (.A(\soc/cpu/_00709_ ),
    .B(\soc/cpu/_02251_ ),
    .Y(\soc/cpu/_04466_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09287_  (.A1(\soc/cpu/reg_next_pc[25] ),
    .A2(net154),
    .B1(\soc/cpu/_04466_ ),
    .Y(\soc/cpu/_04467_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09288_  (.A(\soc/cpu/_04467_ ),
    .Y(\soc/cpu/_04468_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09289_  (.A(\soc/cpu/_04457_ ),
    .B(\soc/cpu/_04468_ ),
    .Y(\soc/cpu/_04469_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09290_  (.A(\soc/cpu/_04443_ ),
    .B(\soc/cpu/_04455_ ),
    .Y(\soc/cpu/_04470_ ));
 sky130_fd_sc_hd__o41a_1 \soc/cpu/_09291_  (.A1(\soc/cpu/_04407_ ),
    .A2(\soc/cpu/_04420_ ),
    .A3(\soc/cpu/_04435_ ),
    .A4(\soc/cpu/_04452_ ),
    .B1(\soc/cpu/decoded_imm_j[20] ),
    .X(\soc/cpu/_04471_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/cpu/_09292_  (.A1(\soc/cpu/_04412_ ),
    .A2(\soc/cpu/_04424_ ),
    .A3(\soc/cpu/_04470_ ),
    .B1(\soc/cpu/_04471_ ),
    .Y(\soc/cpu/_04472_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09293_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04467_ ),
    .Y(\soc/cpu/_04473_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09294_  (.A(\soc/cpu/_04472_ ),
    .B(\soc/cpu/_04473_ ),
    .X(\soc/cpu/_04474_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09295_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04474_ ),
    .B1(\soc/cpu/_03993_ ),
    .Y(\soc/cpu/_04475_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09296_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04469_ ),
    .B1(\soc/cpu/_04475_ ),
    .Y(\soc/cpu/_04476_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09297_  (.A1(\soc/cpu/_04131_ ),
    .A2(\soc/cpu/_04468_ ),
    .B1(\soc/cpu/_04469_ ),
    .B2(\soc/cpu/_03311_ ),
    .Y(\soc/cpu/_04477_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09298_  (.A1(\soc/cpu/_04476_ ),
    .A2(\soc/cpu/_04477_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04478_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09299_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[25] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04468_ ),
    .C1(\soc/cpu/_04478_ ),
    .Y(\soc/cpu/_04479_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09300_  (.A(net131),
    .B(\soc/cpu/_04479_ ),
    .Y(\soc/cpu/_00368_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09301_  (.A1(\soc/cpu/reg_next_pc[26] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04480_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09302_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02254_ ),
    .B1(\soc/cpu/_04480_ ),
    .Y(\soc/cpu/_04481_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09303_  (.A(\soc/cpu/_03300_ ),
    .B(\soc/cpu/_04481_ ),
    .Y(\soc/cpu/_04482_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09304_  (.A(\soc/cpu/_04457_ ),
    .B(\soc/cpu/_04467_ ),
    .Y(\soc/cpu/_04483_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09305_  (.A(\soc/cpu/_04483_ ),
    .B(\soc/cpu/_04481_ ),
    .X(\soc/cpu/_04484_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/cpu/_09306_  (.A_N(\soc/cpu/_04472_ ),
    .B(\soc/cpu/_04473_ ),
    .Y(\soc/cpu/_04485_ ));
 sky130_fd_sc_hd__a21boi_0 \soc/cpu/_09307_  (.A1(\soc/cpu/decoded_imm_j[20] ),
    .A2(\soc/cpu/_04468_ ),
    .B1_N(\soc/cpu/_04485_ ),
    .Y(\soc/cpu/_04486_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09308_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04481_ ),
    .Y(\soc/cpu/_04487_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09309_  (.A(\soc/cpu/_04486_ ),
    .B(\soc/cpu/_04487_ ),
    .Y(\soc/cpu/_04488_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09310_  (.A(\soc/cpu/_04481_ ),
    .SLEEP(\soc/cpu/decoder_trigger ),
    .X(\soc/cpu/_04489_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09311_  (.A1(\soc/cpu/_00818_ ),
    .A2(\soc/cpu/_04484_ ),
    .B1(\soc/cpu/_04489_ ),
    .Y(\soc/cpu/_04490_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09312_  (.A1(\soc/cpu/_00926_ ),
    .A2(\soc/cpu/_04488_ ),
    .B1(\soc/cpu/_04490_ ),
    .Y(\soc/cpu/_04491_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09313_  (.A1(\soc/cpu/_03311_ ),
    .A2(\soc/cpu/_04484_ ),
    .B1(\soc/cpu/_04491_ ),
    .B2(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04492_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09314_  (.A1(\soc/cpu/_04482_ ),
    .A2(\soc/cpu/_04492_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04493_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09315_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[26] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04481_ ),
    .C1(\soc/cpu/_04493_ ),
    .Y(\soc/cpu/_04494_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09316_  (.A(net131),
    .B(\soc/cpu/_04494_ ),
    .Y(\soc/cpu/_00369_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09317_  (.A(\soc/cpu/_00709_ ),
    .B(\soc/cpu/_02260_ ),
    .Y(\soc/cpu/_04495_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09318_  (.A1(\soc/cpu/reg_next_pc[27] ),
    .A2(net154),
    .B1(\soc/cpu/_04495_ ),
    .Y(\soc/cpu/_04496_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09319_  (.A(\soc/cpu/_04496_ ),
    .Y(\soc/cpu/_04497_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09320_  (.A(\soc/cpu/_04483_ ),
    .B(\soc/cpu/_04481_ ),
    .Y(\soc/cpu/_04498_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09321_  (.A(\soc/cpu/_04498_ ),
    .B(\soc/cpu/_04497_ ),
    .Y(\soc/cpu/_04499_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09322_  (.A(\soc/cpu/_03311_ ),
    .B(\soc/cpu/_04499_ ),
    .Y(\soc/cpu/_04500_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09323_  (.A(\soc/cpu/_04131_ ),
    .B(\soc/cpu/_04497_ ),
    .Y(\soc/cpu/_04501_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09324_  (.A1(\soc/cpu/_04468_ ),
    .A2(\soc/cpu/_04481_ ),
    .B1(\soc/cpu/decoded_imm_j[20] ),
    .Y(\soc/cpu/_04502_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09325_  (.A1(\soc/cpu/_04485_ ),
    .A2(\soc/cpu/_04487_ ),
    .B1(\soc/cpu/_04502_ ),
    .Y(\soc/cpu/_04503_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09326_  (.A(\soc/cpu/_02484_ ),
    .B(\soc/cpu/_04496_ ),
    .Y(\soc/cpu/_04504_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09327_  (.A(\soc/cpu/_04503_ ),
    .B(\soc/cpu/_04504_ ),
    .X(\soc/cpu/_04505_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09328_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04505_ ),
    .B1(\soc/cpu/_03993_ ),
    .Y(\soc/cpu/_04506_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09329_  (.A1(\soc/cpu/instr_jal ),
    .A2(\soc/cpu/_04499_ ),
    .B1(\soc/cpu/_04506_ ),
    .Y(\soc/cpu/_04507_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09330_  (.A1(\soc/cpu/_04500_ ),
    .A2(\soc/cpu/_04501_ ),
    .A3(\soc/cpu/_04507_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04508_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/cpu/_09331_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[27] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04497_ ),
    .C1(\soc/cpu/_04508_ ),
    .Y(\soc/cpu/_04509_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09332_  (.A(net131),
    .B(\soc/cpu/_04509_ ),
    .Y(\soc/cpu/_00370_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09333_  (.A(\soc/cpu/_01731_ ),
    .B(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04510_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09334_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02263_ ),
    .B1(\soc/cpu/_04510_ ),
    .Y(\soc/cpu/_04511_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09335_  (.A(\soc/cpu/_03300_ ),
    .B(\soc/cpu/_04511_ ),
    .Y(\soc/cpu/_04512_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09336_  (.A(\soc/cpu/_04498_ ),
    .B(\soc/cpu/_04496_ ),
    .Y(\soc/cpu/_04513_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09337_  (.A(\soc/cpu/_04513_ ),
    .B(\soc/cpu/_04511_ ),
    .X(\soc/cpu/_04514_ ));
 sky130_fd_sc_hd__maj3_1 \soc/cpu/_09338_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04503_ ),
    .C(\soc/cpu/_04497_ ),
    .X(\soc/cpu/_04515_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09339_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04511_ ),
    .Y(\soc/cpu/_04516_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09340_  (.A(\soc/cpu/_04515_ ),
    .B(\soc/cpu/_04516_ ),
    .X(\soc/cpu/_04517_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09341_  (.A(\soc/cpu/_04511_ ),
    .SLEEP(\soc/cpu/decoder_trigger ),
    .X(\soc/cpu/_04518_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09342_  (.A1(\soc/cpu/_00818_ ),
    .A2(\soc/cpu/_04514_ ),
    .B1(\soc/cpu/_04518_ ),
    .Y(\soc/cpu/_04519_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09343_  (.A1(\soc/cpu/_00926_ ),
    .A2(\soc/cpu/_04517_ ),
    .B1(\soc/cpu/_04519_ ),
    .Y(\soc/cpu/_04520_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09344_  (.A1(\soc/cpu/_03311_ ),
    .A2(\soc/cpu/_04514_ ),
    .B1(\soc/cpu/_04520_ ),
    .B2(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04521_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09345_  (.A1(\soc/cpu/_04512_ ),
    .A2(\soc/cpu/_04521_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04522_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09346_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[28] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04511_ ),
    .X(\soc/cpu/_04523_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09347_  (.A1(\soc/cpu/_04522_ ),
    .A2(\soc/cpu/_04523_ ),
    .B1(_074_),
    .X(\soc/cpu/_00371_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09348_  (.A(\soc/cpu/_04504_ ),
    .B(\soc/cpu/_04516_ ),
    .Y(\soc/cpu/_04524_ ));
 sky130_fd_sc_hd__nor4bb_1 \soc/cpu/_09349_  (.A(\soc/cpu/_04487_ ),
    .B(\soc/cpu/_04472_ ),
    .C_N(\soc/cpu/_04473_ ),
    .D_N(\soc/cpu/_04524_ ),
    .Y(\soc/cpu/_04525_ ));
 sky130_fd_sc_hd__o41a_1 \soc/cpu/_09350_  (.A1(\soc/cpu/_04468_ ),
    .A2(\soc/cpu/_04481_ ),
    .A3(\soc/cpu/_04497_ ),
    .A4(\soc/cpu/_04511_ ),
    .B1(\soc/cpu/decoded_imm_j[20] ),
    .X(\soc/cpu/_04526_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09351_  (.A(\soc/cpu/_00709_ ),
    .B(\soc/cpu/_02269_ ),
    .Y(\soc/cpu/_04527_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09352_  (.A1(\soc/cpu/reg_next_pc[29] ),
    .A2(\soc/cpu/_04116_ ),
    .B1(\soc/cpu/_04527_ ),
    .Y(\soc/cpu/_04528_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09353_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04528_ ),
    .Y(\soc/cpu/_04529_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09354_  (.A1(\soc/cpu/_04525_ ),
    .A2(\soc/cpu/_04526_ ),
    .B1(\soc/cpu/_04529_ ),
    .Y(\soc/cpu/_04530_ ));
 sky130_fd_sc_hd__or3_1 \soc/cpu/_09355_  (.A(\soc/cpu/_04525_ ),
    .B(\soc/cpu/_04526_ ),
    .C(\soc/cpu/_04529_ ),
    .X(\soc/cpu/_04531_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09356_  (.A(\soc/cpu/_03312_ ),
    .B(\soc/cpu/_04530_ ),
    .C(\soc/cpu/_04531_ ),
    .Y(\soc/cpu/_04532_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09357_  (.A(\soc/cpu/_04513_ ),
    .B(\soc/cpu/_04511_ ),
    .Y(\soc/cpu/_04533_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09358_  (.A(\soc/cpu/_04533_ ),
    .B(\soc/cpu/_04528_ ),
    .X(\soc/cpu/_04534_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09359_  (.A(\soc/cpu/_03311_ ),
    .B(\soc/cpu/_04534_ ),
    .Y(\soc/cpu/_04535_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09360_  (.A(\soc/cpu/_00928_ ),
    .B(\soc/cpu/_03311_ ),
    .C(\soc/cpu/_04528_ ),
    .Y(\soc/cpu/_04536_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09361_  (.A1(\soc/cpu/_03323_ ),
    .A2(\soc/cpu/_04534_ ),
    .B1(\soc/cpu/_04536_ ),
    .Y(\soc/cpu/_04537_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09362_  (.A1(\soc/cpu/_04532_ ),
    .A2(\soc/cpu/_04535_ ),
    .A3(\soc/cpu/_04537_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04538_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09363_  (.A(\soc/cpu/_00953_ ),
    .B(\soc/cpu/_04528_ ),
    .Y(\soc/cpu/_04539_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_09364_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[29] ),
    .B1(\soc/cpu/_04538_ ),
    .C1(\soc/cpu/_04539_ ),
    .Y(\soc/cpu/_04540_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09365_  (.A(net132),
    .B(\soc/cpu/_04540_ ),
    .Y(\soc/cpu/_00372_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09366_  (.A(\soc/cpu/_00709_ ),
    .B(\soc/cpu/_02274_ ),
    .Y(\soc/cpu/_04541_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/_09367_  (.A1(\soc/cpu/reg_next_pc[30] ),
    .A2(\soc/cpu/_04116_ ),
    .B1(\soc/cpu/_04541_ ),
    .Y(\soc/cpu/_04542_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09368_  (.A(\soc/cpu/_04542_ ),
    .Y(\soc/cpu/_04543_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09369_  (.A(\soc/cpu/_03300_ ),
    .B(\soc/cpu/_04543_ ),
    .Y(\soc/cpu/_04544_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09370_  (.A(\soc/cpu/_04533_ ),
    .B(\soc/cpu/_04528_ ),
    .Y(\soc/cpu/_04545_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09371_  (.A(\soc/cpu/_04545_ ),
    .B(\soc/cpu/_04542_ ),
    .Y(\soc/cpu/_04546_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09372_  (.A1(\soc/cpu/_02484_ ),
    .A2(\soc/cpu/_04528_ ),
    .B1(\soc/cpu/_04530_ ),
    .Y(\soc/cpu/_04547_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09373_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04542_ ),
    .Y(\soc/cpu/_04548_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09374_  (.A(\soc/cpu/_04547_ ),
    .B(\soc/cpu/_04548_ ),
    .Y(\soc/cpu/_04549_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09375_  (.A(\soc/cpu/_00818_ ),
    .B(\soc/cpu/_04546_ ),
    .Y(\soc/cpu/_04550_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/_09376_  (.A1(\soc/cpu/decoder_trigger ),
    .A2(\soc/cpu/_04542_ ),
    .B1(\soc/cpu/_04549_ ),
    .B2(\soc/cpu/_00926_ ),
    .C1(\soc/cpu/_04550_ ),
    .Y(\soc/cpu/_04551_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09377_  (.A1(\soc/cpu/_03311_ ),
    .A2(\soc/cpu/_04546_ ),
    .B1(\soc/cpu/_04551_ ),
    .B2(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04552_ ));
 sky130_fd_sc_hd__a21o_1 \soc/cpu/_09378_  (.A1(\soc/cpu/_04544_ ),
    .A2(\soc/cpu/_04552_ ),
    .B1(\soc/cpu/_03994_ ),
    .X(\soc/cpu/_04553_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09379_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[30] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04543_ ),
    .Y(\soc/cpu/_04554_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09380_  (.A1(\soc/cpu/_04553_ ),
    .A2(\soc/cpu/_04554_ ),
    .B1(net131),
    .Y(\soc/cpu/_00373_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09381_  (.A(\soc/cpu/decoded_imm_j[20] ),
    .B(\soc/cpu/_04543_ ),
    .Y(\soc/cpu/_04555_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09382_  (.A1(\soc/cpu/reg_next_pc[31] ),
    .A2(\soc/cpu/_00707_ ),
    .B1(\soc/cpu/_04136_ ),
    .Y(\soc/cpu/_04556_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/cpu/_09383_  (.A1(\soc/cpu/_00707_ ),
    .A2(\soc/cpu/_02279_ ),
    .B1(\soc/cpu/_04556_ ),
    .Y(\soc/cpu/_04557_ ));
 sky130_fd_sc_hd__or4b_1 \soc/cpu/_09384_  (.A(\soc/cpu/_02484_ ),
    .B(\soc/cpu/_04525_ ),
    .C(\soc/cpu/_04526_ ),
    .D_N(\soc/cpu/_04528_ ),
    .X(\soc/cpu/_04558_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/_09385_  (.A1(\soc/cpu/_04530_ ),
    .A2(\soc/cpu/_04542_ ),
    .B1(\soc/cpu/_04558_ ),
    .Y(\soc/cpu/_04559_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09386_  (.A(\soc/cpu/_04555_ ),
    .B(\soc/cpu/_04557_ ),
    .C(\soc/cpu/_04559_ ),
    .X(\soc/cpu/_04560_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09387_  (.A1(\soc/cpu/_04555_ ),
    .A2(\soc/cpu/_04559_ ),
    .B1(\soc/cpu/_04557_ ),
    .Y(\soc/cpu/_04561_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09388_  (.A(\soc/cpu/_00926_ ),
    .B(\soc/cpu/_04560_ ),
    .C(\soc/cpu/_04561_ ),
    .Y(\soc/cpu/_04562_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09389_  (.A(\soc/cpu/_04557_ ),
    .Y(\soc/cpu/_04563_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09390_  (.A(\soc/cpu/_04545_ ),
    .B(\soc/cpu/_04543_ ),
    .Y(\soc/cpu/_04564_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09391_  (.A(\soc/cpu/_04564_ ),
    .B(\soc/cpu/_04563_ ),
    .Y(\soc/cpu/_04565_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/_09392_  (.A1(\soc/cpu/decoder_trigger ),
    .A2(\soc/cpu/_04563_ ),
    .B1(\soc/cpu/_04565_ ),
    .B2(\soc/cpu/_03322_ ),
    .Y(\soc/cpu/_04566_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09393_  (.A1(\soc/cpu/_04562_ ),
    .A2(\soc/cpu/_04566_ ),
    .B1(\soc/cpu/_00797_ ),
    .Y(\soc/cpu/_04567_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09394_  (.A(\soc/cpu/_03403_ ),
    .B(\soc/cpu/_04565_ ),
    .Y(\soc/cpu/_04568_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09395_  (.A1(\soc/cpu/_03300_ ),
    .A2(\soc/cpu/_04557_ ),
    .B1(\soc/cpu/_04568_ ),
    .Y(\soc/cpu/_04569_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09396_  (.A1(\soc/cpu/_04567_ ),
    .A2(\soc/cpu/_04569_ ),
    .B1(\soc/cpu/_03994_ ),
    .Y(\soc/cpu/_04570_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09397_  (.A1(\soc/cpu/_00839_ ),
    .A2(\soc/cpu/reg_next_pc[31] ),
    .B1(\soc/cpu/_04114_ ),
    .B2(\soc/cpu/_04557_ ),
    .X(\soc/cpu/_04571_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09398_  (.A1(\soc/cpu/_04570_ ),
    .A2(\soc/cpu/_04571_ ),
    .B1(_074_),
    .X(\soc/cpu/_00374_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09401_  (.A(\soc/cpu/reg_pc[1] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04574_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09402_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04122_ ),
    .B1(\soc/cpu/_04574_ ),
    .Y(\soc/cpu/_00375_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09403_  (.A(\soc/cpu/reg_pc[2] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04575_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09404_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04133_ ),
    .B1(\soc/cpu/_04575_ ),
    .Y(\soc/cpu/_00376_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09405_  (.A(\soc/cpu/reg_pc[3] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04576_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09406_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04146_ ),
    .B1(\soc/cpu/_04576_ ),
    .Y(\soc/cpu/_00377_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09408_  (.A1(\soc/cpu/reg_pc[4] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04162_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00378_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09409_  (.A1(\soc/cpu/reg_pc[5] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04172_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00379_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09410_  (.A1(\soc/cpu/reg_pc[6] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04184_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00380_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09411_  (.A1(\soc/cpu/reg_pc[7] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04195_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00381_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09412_  (.A1(\soc/cpu/reg_pc[8] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04209_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00382_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09413_  (.A1(\soc/cpu/reg_pc[9] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04226_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00383_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09414_  (.A1(\soc/cpu/reg_pc[10] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04241_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00384_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09415_  (.A1(\soc/cpu/reg_pc[11] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04254_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00385_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09417_  (.A1(\soc/cpu/reg_pc[12] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04267_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00386_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09418_  (.A1(\soc/cpu/reg_pc[13] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04284_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00387_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09419_  (.A(\soc/cpu/reg_pc[14] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04579_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09420_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04306_ ),
    .B1(\soc/cpu/_04579_ ),
    .Y(\soc/cpu/_00388_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09422_  (.A1(\soc/cpu/reg_pc[15] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04316_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00389_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09423_  (.A1(\soc/cpu/reg_pc[16] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04332_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00390_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09424_  (.A1(\soc/cpu/reg_pc[17] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04349_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00391_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09425_  (.A(\soc/cpu/reg_pc[18] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04581_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09426_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04367_ ),
    .B1(\soc/cpu/_04581_ ),
    .Y(\soc/cpu/_00392_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09427_  (.A1(\soc/cpu/reg_pc[19] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04377_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00393_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09428_  (.A1(\soc/cpu/reg_pc[20] ),
    .A2(\soc/cpu/_03330_ ),
    .B1(\soc/cpu/_04390_ ),
    .B2(\soc/cpu/_00795_ ),
    .X(\soc/cpu/_00394_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09429_  (.A1(\soc/cpu/reg_pc[21] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04407_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00395_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09430_  (.A1(\soc/cpu/reg_pc[22] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04420_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00396_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09431_  (.A1(\soc/cpu/reg_pc[23] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04435_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00397_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09432_  (.A1(\soc/cpu/reg_pc[24] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04452_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00398_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09433_  (.A(\soc/cpu/reg_pc[25] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04582_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09434_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04467_ ),
    .B1(\soc/cpu/_04582_ ),
    .Y(\soc/cpu/_00399_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09435_  (.A1(\soc/cpu/reg_pc[26] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04481_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00400_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09436_  (.A(\soc/cpu/reg_pc[27] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04583_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09437_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04496_ ),
    .B1(\soc/cpu/_04583_ ),
    .Y(\soc/cpu/_00401_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/_09438_  (.A1(\soc/cpu/reg_pc[28] ),
    .A2(\soc/cpu/_03303_ ),
    .B1(\soc/cpu/_04511_ ),
    .B2(\soc/cpu/_00859_ ),
    .X(\soc/cpu/_00402_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09439_  (.A(\soc/cpu/reg_pc[29] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04584_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09440_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04528_ ),
    .B1(\soc/cpu/_04584_ ),
    .Y(\soc/cpu/_00403_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09441_  (.A(\soc/cpu/reg_pc[30] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04585_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09442_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04542_ ),
    .B1(\soc/cpu/_04585_ ),
    .Y(\soc/cpu/_00404_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09443_  (.A(\soc/cpu/reg_pc[31] ),
    .B(\soc/cpu/_03303_ ),
    .Y(\soc/cpu/_04586_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09444_  (.A1(\soc/cpu/_00795_ ),
    .A2(\soc/cpu/_04563_ ),
    .B1(\soc/cpu/_04586_ ),
    .Y(\soc/cpu/_00405_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09445_  (.A1(\soc/cpu/count_instr[0] ),
    .A2(\soc/cpu/_03995_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04587_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09446_  (.A1(\soc/cpu/count_instr[0] ),
    .A2(\soc/cpu/_03995_ ),
    .B1(\soc/cpu/_04587_ ),
    .Y(\soc/cpu/_00406_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09448_  (.A(\soc/cpu/count_instr[0] ),
    .B(\soc/cpu/count_instr[1] ),
    .C(\soc/cpu/_03995_ ),
    .X(\soc/cpu/_04589_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09449_  (.A1(\soc/cpu/count_instr[0] ),
    .A2(\soc/cpu/_03995_ ),
    .B1(\soc/cpu/count_instr[1] ),
    .Y(\soc/cpu/_04590_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09450_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04589_ ),
    .C(\soc/cpu/_04590_ ),
    .Y(\soc/cpu/_00407_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09451_  (.A(\soc/cpu/count_instr[2] ),
    .B(\soc/cpu/_04589_ ),
    .X(\soc/cpu/_04591_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09452_  (.A1(\soc/cpu/count_instr[2] ),
    .A2(\soc/cpu/_04589_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04592_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09453_  (.A(\soc/cpu/_04591_ ),
    .B(\soc/cpu/_04592_ ),
    .Y(\soc/cpu/_00408_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09454_  (.A1(\soc/cpu/count_instr[3] ),
    .A2(\soc/cpu/_04591_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04593_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09455_  (.A(\soc/cpu/count_instr[2] ),
    .B(\soc/cpu/count_instr[3] ),
    .C(\soc/cpu/_04589_ ),
    .X(\soc/cpu/_04594_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09456_  (.A(\soc/cpu/_04593_ ),
    .B(\soc/cpu/_04594_ ),
    .Y(\soc/cpu/_00409_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09457_  (.A1(\soc/cpu/count_instr[4] ),
    .A2(\soc/cpu/_04594_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04595_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09458_  (.A(\soc/cpu/count_instr[3] ),
    .B(\soc/cpu/count_instr[4] ),
    .C(\soc/cpu/_04591_ ),
    .X(\soc/cpu/_04596_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09459_  (.A(\soc/cpu/_04595_ ),
    .B(\soc/cpu/_04596_ ),
    .Y(\soc/cpu/_00410_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09460_  (.A1(\soc/cpu/count_instr[5] ),
    .A2(\soc/cpu/_04596_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04597_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09461_  (.A1(\soc/cpu/count_instr[5] ),
    .A2(\soc/cpu/_04596_ ),
    .B1(\soc/cpu/_04597_ ),
    .Y(\soc/cpu/_00411_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09462_  (.A1(\soc/cpu/count_instr[5] ),
    .A2(\soc/cpu/_04596_ ),
    .B1(\soc/cpu/count_instr[6] ),
    .Y(\soc/cpu/_04598_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09463_  (.A(\soc/cpu/count_instr[4] ),
    .B(\soc/cpu/_04594_ ),
    .Y(\soc/cpu/_04599_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09464_  (.A(\soc/cpu/count_instr[5] ),
    .B(\soc/cpu/count_instr[6] ),
    .Y(\soc/cpu/_04600_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09465_  (.A(\soc/cpu/_04599_ ),
    .B(\soc/cpu/_04600_ ),
    .Y(\soc/cpu/_04601_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09466_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04598_ ),
    .C(\soc/cpu/_04601_ ),
    .Y(\soc/cpu/_00412_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09467_  (.A1(\soc/cpu/count_instr[7] ),
    .A2(\soc/cpu/_04601_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04602_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09468_  (.A(\soc/cpu/count_instr[7] ),
    .B(\soc/cpu/_04601_ ),
    .X(\soc/cpu/_04603_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09469_  (.A(\soc/cpu/_04602_ ),
    .B(\soc/cpu/_04603_ ),
    .Y(\soc/cpu/_00413_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09470_  (.A1(\soc/cpu/count_instr[8] ),
    .A2(\soc/cpu/_04603_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04604_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09471_  (.A(\soc/cpu/count_instr[7] ),
    .B(\soc/cpu/count_instr[8] ),
    .C(\soc/cpu/_04601_ ),
    .X(\soc/cpu/_04605_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09472_  (.A(\soc/cpu/_04604_ ),
    .B(\soc/cpu/_04605_ ),
    .Y(\soc/cpu/_00414_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09473_  (.A1(\soc/cpu/count_instr[9] ),
    .A2(\soc/cpu/_04605_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04606_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09474_  (.A(\soc/cpu/count_instr[8] ),
    .B(\soc/cpu/count_instr[9] ),
    .C(\soc/cpu/_04603_ ),
    .X(\soc/cpu/_04607_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09475_  (.A(\soc/cpu/_04606_ ),
    .B(\soc/cpu/_04607_ ),
    .Y(\soc/cpu/_00415_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09476_  (.A1(\soc/cpu/count_instr[10] ),
    .A2(\soc/cpu/_04607_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04608_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09477_  (.A1(\soc/cpu/count_instr[10] ),
    .A2(\soc/cpu/_04607_ ),
    .B1(\soc/cpu/_04608_ ),
    .Y(\soc/cpu/_00416_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09478_  (.A(\soc/cpu/count_instr[1] ),
    .B(\soc/cpu/count_instr[2] ),
    .C(\soc/cpu/count_instr[4] ),
    .X(\soc/cpu/_04609_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09479_  (.A(\soc/cpu/count_instr[0] ),
    .B(\soc/cpu/count_instr[3] ),
    .C(\soc/cpu/_03995_ ),
    .D(\soc/cpu/_04609_ ),
    .Y(\soc/cpu/_04610_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09480_  (.A(\soc/cpu/count_instr[7] ),
    .B(\soc/cpu/count_instr[8] ),
    .C(\soc/cpu/count_instr[9] ),
    .D(\soc/cpu/count_instr[10] ),
    .Y(\soc/cpu/_04611_ ));
 sky130_fd_sc_hd__or2_2 \soc/cpu/_09481_  (.A(\soc/cpu/_04600_ ),
    .B(\soc/cpu/_04611_ ),
    .X(\soc/cpu/_04612_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09482_  (.A(\soc/cpu/_04610_ ),
    .B(\soc/cpu/_04612_ ),
    .Y(\soc/cpu/_04613_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09483_  (.A1(\soc/cpu/count_instr[11] ),
    .A2(\soc/cpu/_04613_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04614_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09484_  (.A1(\soc/cpu/count_instr[11] ),
    .A2(\soc/cpu/_04613_ ),
    .B1(\soc/cpu/_04614_ ),
    .Y(\soc/cpu/_00417_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09485_  (.A1(\soc/cpu/count_instr[11] ),
    .A2(\soc/cpu/_04613_ ),
    .B1(\soc/cpu/count_instr[12] ),
    .Y(\soc/cpu/_04615_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09486_  (.A(\soc/cpu/count_instr[11] ),
    .B(net785),
    .Y(\soc/cpu/_04616_ ));
 sky130_fd_sc_hd__nor3_2 \soc/cpu/_09487_  (.A(\soc/cpu/_04599_ ),
    .B(\soc/cpu/_04612_ ),
    .C(net786),
    .Y(\soc/cpu/_04617_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09488_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04615_ ),
    .C(\soc/cpu/_04617_ ),
    .Y(\soc/cpu/_00418_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09489_  (.A1(\soc/cpu/count_instr[13] ),
    .A2(\soc/cpu/_04617_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04618_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09490_  (.A1(\soc/cpu/count_instr[13] ),
    .A2(\soc/cpu/_04617_ ),
    .B1(\soc/cpu/_04618_ ),
    .Y(\soc/cpu/_00419_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09491_  (.A1(net760),
    .A2(\soc/cpu/_04617_ ),
    .B1(\soc/cpu/count_instr[14] ),
    .Y(\soc/cpu/_04619_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09492_  (.A(net760),
    .B(\soc/cpu/count_instr[14] ),
    .C(\soc/cpu/_04617_ ),
    .X(\soc/cpu/_04620_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09493_  (.A(\soc/cpu/_00840_ ),
    .B(net761),
    .C(\soc/cpu/_04620_ ),
    .Y(\soc/cpu/_00420_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09494_  (.A1(\soc/cpu/count_instr[15] ),
    .A2(\soc/cpu/_04620_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04621_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09495_  (.A1(\soc/cpu/count_instr[15] ),
    .A2(\soc/cpu/_04620_ ),
    .B1(\soc/cpu/_04621_ ),
    .Y(\soc/cpu/_00421_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09496_  (.A(net798),
    .B(net785),
    .C(\soc/cpu/_04613_ ),
    .Y(\soc/cpu/_04622_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09497_  (.A(net760),
    .B(\soc/cpu/count_instr[14] ),
    .C(\soc/cpu/count_instr[15] ),
    .Y(\soc/cpu/_04623_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09498_  (.A(\soc/cpu/_04622_ ),
    .B(\soc/cpu/_04623_ ),
    .Y(\soc/cpu/_04624_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09499_  (.A1(\soc/cpu/count_instr[16] ),
    .A2(\soc/cpu/_04624_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04625_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09500_  (.A1(\soc/cpu/count_instr[16] ),
    .A2(\soc/cpu/_04624_ ),
    .B1(\soc/cpu/_04625_ ),
    .Y(\soc/cpu/_00422_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09501_  (.A1(\soc/cpu/count_instr[16] ),
    .A2(\soc/cpu/_04624_ ),
    .B1(\soc/cpu/count_instr[17] ),
    .Y(\soc/cpu/_04626_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09502_  (.A(\soc/cpu/count_instr[16] ),
    .B(\soc/cpu/count_instr[17] ),
    .C(\soc/cpu/_04624_ ),
    .X(\soc/cpu/_04627_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09503_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04626_ ),
    .C(\soc/cpu/_04627_ ),
    .Y(\soc/cpu/_00423_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09505_  (.A1(\soc/cpu/count_instr[18] ),
    .A2(\soc/cpu/_04627_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04629_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09506_  (.A(\soc/cpu/count_instr[18] ),
    .B(\soc/cpu/_04627_ ),
    .X(\soc/cpu/_04630_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09507_  (.A(\soc/cpu/_04629_ ),
    .B(\soc/cpu/_04630_ ),
    .Y(\soc/cpu/_00424_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09508_  (.A1(\soc/cpu/count_instr[19] ),
    .A2(\soc/cpu/_04630_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04631_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09509_  (.A1(\soc/cpu/count_instr[19] ),
    .A2(\soc/cpu/_04630_ ),
    .B1(\soc/cpu/_04631_ ),
    .Y(\soc/cpu/_00425_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09510_  (.A(\soc/cpu/count_instr[16] ),
    .B(\soc/cpu/count_instr[17] ),
    .C(\soc/cpu/count_instr[18] ),
    .D(\soc/cpu/count_instr[19] ),
    .Y(\soc/cpu/_04632_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09511_  (.A(net786),
    .B(\soc/cpu/_04623_ ),
    .C(\soc/cpu/_04632_ ),
    .Y(\soc/cpu/_04633_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09512_  (.A1(\soc/cpu/_04613_ ),
    .A2(\soc/cpu/_04633_ ),
    .B1(\soc/cpu/count_instr[20] ),
    .Y(\soc/cpu/_04634_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09513_  (.A(\soc/cpu/_04599_ ),
    .B(\soc/cpu/_04612_ ),
    .Y(\soc/cpu/_04635_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09514_  (.A(\soc/cpu/count_instr[20] ),
    .B(\soc/cpu/_04635_ ),
    .C(\soc/cpu/_04633_ ),
    .X(\soc/cpu/_04636_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09515_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04634_ ),
    .C(\soc/cpu/_04636_ ),
    .Y(\soc/cpu/_00426_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09516_  (.A1(\soc/cpu/count_instr[21] ),
    .A2(\soc/cpu/_04636_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04637_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09517_  (.A1(\soc/cpu/count_instr[21] ),
    .A2(\soc/cpu/_04636_ ),
    .B1(\soc/cpu/_04637_ ),
    .Y(\soc/cpu/_00427_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09518_  (.A1(\soc/cpu/count_instr[21] ),
    .A2(\soc/cpu/_04636_ ),
    .B1(\soc/cpu/count_instr[22] ),
    .Y(\soc/cpu/_04638_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09519_  (.A(\soc/cpu/count_instr[21] ),
    .B(\soc/cpu/count_instr[22] ),
    .C(\soc/cpu/_04636_ ),
    .X(\soc/cpu/_04639_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09520_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04638_ ),
    .C(\soc/cpu/_04639_ ),
    .Y(\soc/cpu/_00428_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09521_  (.A1(\soc/cpu/count_instr[23] ),
    .A2(\soc/cpu/_04639_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04640_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09522_  (.A(\soc/cpu/count_instr[23] ),
    .B(\soc/cpu/_04639_ ),
    .X(\soc/cpu/_04641_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09523_  (.A(\soc/cpu/_04640_ ),
    .B(\soc/cpu/_04641_ ),
    .Y(\soc/cpu/_00429_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09524_  (.A1(\soc/cpu/count_instr[24] ),
    .A2(\soc/cpu/_04641_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04642_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09525_  (.A1(\soc/cpu/count_instr[23] ),
    .A2(\soc/cpu/count_instr[24] ),
    .A3(\soc/cpu/_04639_ ),
    .B1(\soc/cpu/_04642_ ),
    .Y(\soc/cpu/_00430_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09526_  (.A(\soc/cpu/count_instr[23] ),
    .B(\soc/cpu/count_instr[24] ),
    .C(\soc/cpu/count_instr[25] ),
    .Y(\soc/cpu/_04643_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09527_  (.A(\soc/cpu/count_instr[0] ),
    .B(\soc/cpu/count_instr[1] ),
    .C(\soc/cpu/count_instr[4] ),
    .Y(\soc/cpu/_04644_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09528_  (.A(\soc/cpu/count_instr[2] ),
    .B(\soc/cpu/count_instr[3] ),
    .C(\soc/cpu/count_instr[21] ),
    .D(\soc/cpu/count_instr[22] ),
    .Y(\soc/cpu/_04645_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_09529_  (.A(\soc/cpu/_04612_ ),
    .B(\soc/cpu/_04643_ ),
    .C(\soc/cpu/_04644_ ),
    .D(\soc/cpu/_04645_ ),
    .Y(\soc/cpu/_04646_ ));
 sky130_fd_sc_hd__nand3_2 \soc/cpu/_09530_  (.A(\soc/cpu/count_instr[20] ),
    .B(\soc/cpu/_04633_ ),
    .C(\soc/cpu/_04646_ ),
    .Y(\soc/cpu/_04647_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/_09531_  (.A(\soc/cpu/_03993_ ),
    .B(\soc/cpu/_03994_ ),
    .C(\soc/cpu/_04647_ ),
    .Y(\soc/cpu/_04648_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09532_  (.A1(\soc/cpu/count_instr[23] ),
    .A2(\soc/cpu/count_instr[24] ),
    .A3(\soc/cpu/_04639_ ),
    .B1(\soc/cpu/count_instr[25] ),
    .Y(\soc/cpu/_04649_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09533_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04648_ ),
    .C(\soc/cpu/_04649_ ),
    .Y(\soc/cpu/_00431_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09534_  (.A1(\soc/cpu/count_instr[26] ),
    .A2(\soc/cpu/_04648_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04650_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09535_  (.A1(\soc/cpu/count_instr[26] ),
    .A2(\soc/cpu/_04648_ ),
    .B1(\soc/cpu/_04650_ ),
    .Y(\soc/cpu/_00432_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09536_  (.A1(\soc/cpu/count_instr[26] ),
    .A2(\soc/cpu/_04648_ ),
    .B1(\soc/cpu/count_instr[27] ),
    .Y(\soc/cpu/_04651_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09537_  (.A(\soc/cpu/count_instr[26] ),
    .B(\soc/cpu/count_instr[27] ),
    .C(\soc/cpu/_04648_ ),
    .X(\soc/cpu/_04652_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09538_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04651_ ),
    .C(\soc/cpu/_04652_ ),
    .Y(\soc/cpu/_00433_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09539_  (.A1(\soc/cpu/count_instr[28] ),
    .A2(\soc/cpu/_04652_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04653_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09540_  (.A(\soc/cpu/count_instr[26] ),
    .B(\soc/cpu/count_instr[27] ),
    .C(\soc/cpu/count_instr[28] ),
    .D(\soc/cpu/_04648_ ),
    .X(\soc/cpu/_04654_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09541_  (.A(\soc/cpu/_04653_ ),
    .B(\soc/cpu/_04654_ ),
    .Y(\soc/cpu/_00434_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09542_  (.A1(\soc/cpu/count_instr[29] ),
    .A2(\soc/cpu/_04654_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04655_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09543_  (.A(\soc/cpu/count_instr[28] ),
    .B(\soc/cpu/count_instr[29] ),
    .C(\soc/cpu/_04652_ ),
    .X(\soc/cpu/_04656_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09544_  (.A(\soc/cpu/_04655_ ),
    .B(\soc/cpu/_04656_ ),
    .Y(\soc/cpu/_00435_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09545_  (.A1(\soc/cpu/count_instr[30] ),
    .A2(\soc/cpu/_04656_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04657_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09546_  (.A(\soc/cpu/count_instr[30] ),
    .B(\soc/cpu/_04656_ ),
    .X(\soc/cpu/_04658_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09547_  (.A(\soc/cpu/_04657_ ),
    .B(\soc/cpu/_04658_ ),
    .Y(\soc/cpu/_00436_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09548_  (.A1(\soc/cpu/count_instr[31] ),
    .A2(\soc/cpu/_04658_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04659_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09549_  (.A(\soc/cpu/count_instr[30] ),
    .B(\soc/cpu/count_instr[31] ),
    .C(\soc/cpu/_04656_ ),
    .X(\soc/cpu/_04660_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09550_  (.A(\soc/cpu/_04659_ ),
    .B(\soc/cpu/_04660_ ),
    .Y(\soc/cpu/_00437_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09551_  (.A1(\soc/cpu/count_instr[32] ),
    .A2(\soc/cpu/_04660_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04661_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09552_  (.A(\soc/cpu/count_instr[29] ),
    .B(\soc/cpu/count_instr[30] ),
    .C(\soc/cpu/count_instr[31] ),
    .X(\soc/cpu/_04662_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09553_  (.A(\soc/cpu/count_instr[32] ),
    .B(\soc/cpu/count_instr[28] ),
    .C(\soc/cpu/_04652_ ),
    .D(\soc/cpu/_04662_ ),
    .X(\soc/cpu/_04663_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09554_  (.A(\soc/cpu/_04661_ ),
    .B(\soc/cpu/_04663_ ),
    .Y(\soc/cpu/_00438_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09555_  (.A1(\soc/cpu/count_instr[33] ),
    .A2(\soc/cpu/_04663_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04664_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09556_  (.A(\soc/cpu/count_instr[32] ),
    .B(\soc/cpu/count_instr[33] ),
    .C(\soc/cpu/_04660_ ),
    .X(\soc/cpu/_04665_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09557_  (.A(\soc/cpu/_04664_ ),
    .B(\soc/cpu/_04665_ ),
    .Y(\soc/cpu/_00439_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09558_  (.A1(\soc/cpu/count_instr[34] ),
    .A2(\soc/cpu/_04665_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04666_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09559_  (.A(\soc/cpu/count_instr[33] ),
    .B(\soc/cpu/count_instr[34] ),
    .C(\soc/cpu/_04663_ ),
    .X(\soc/cpu/_04667_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09560_  (.A(\soc/cpu/_04666_ ),
    .B(\soc/cpu/_04667_ ),
    .Y(\soc/cpu/_00440_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09561_  (.A1(\soc/cpu/count_instr[35] ),
    .A2(\soc/cpu/_04667_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04668_ ));
 sky130_fd_sc_hd__and2_2 \soc/cpu/_09562_  (.A(\soc/cpu/count_instr[35] ),
    .B(\soc/cpu/_04667_ ),
    .X(\soc/cpu/_04669_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09563_  (.A(\soc/cpu/_04668_ ),
    .B(\soc/cpu/_04669_ ),
    .Y(\soc/cpu/_00441_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09565_  (.A1(\soc/cpu/count_instr[36] ),
    .A2(\soc/cpu/_04669_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04671_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09566_  (.A(\soc/cpu/count_instr[35] ),
    .B(\soc/cpu/count_instr[36] ),
    .C(\soc/cpu/_04667_ ),
    .X(\soc/cpu/_04672_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09567_  (.A(\soc/cpu/_04671_ ),
    .B(\soc/cpu/_04672_ ),
    .Y(\soc/cpu/_00442_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09568_  (.A1(\soc/cpu/count_instr[37] ),
    .A2(\soc/cpu/_04672_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04673_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09569_  (.A1(\soc/cpu/count_instr[37] ),
    .A2(\soc/cpu/_04672_ ),
    .B1(\soc/cpu/_04673_ ),
    .Y(\soc/cpu/_00443_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09570_  (.A1(\soc/cpu/count_instr[37] ),
    .A2(\soc/cpu/_04672_ ),
    .B1(\soc/cpu/count_instr[38] ),
    .Y(\soc/cpu/_04674_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09571_  (.A(\soc/cpu/count_instr[36] ),
    .B(\soc/cpu/count_instr[37] ),
    .C(\soc/cpu/count_instr[38] ),
    .D(\soc/cpu/_04669_ ),
    .X(\soc/cpu/_04675_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09572_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04674_ ),
    .C(\soc/cpu/_04675_ ),
    .Y(\soc/cpu/_00444_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09573_  (.A1(\soc/cpu/count_instr[39] ),
    .A2(\soc/cpu/_04675_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04676_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09574_  (.A1(\soc/cpu/count_instr[39] ),
    .A2(\soc/cpu/_04675_ ),
    .B1(\soc/cpu/_04676_ ),
    .Y(\soc/cpu/_00445_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09575_  (.A1(\soc/cpu/count_instr[39] ),
    .A2(\soc/cpu/_04675_ ),
    .B1(\soc/cpu/count_instr[40] ),
    .Y(\soc/cpu/_04677_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09576_  (.A(\soc/cpu/count_instr[36] ),
    .B(\soc/cpu/count_instr[37] ),
    .C(\soc/cpu/count_instr[38] ),
    .D(\soc/cpu/_04669_ ),
    .Y(\soc/cpu/_04678_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09577_  (.A(\soc/cpu/count_instr[39] ),
    .B(\soc/cpu/count_instr[40] ),
    .Y(\soc/cpu/_04679_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09578_  (.A(\soc/cpu/_04678_ ),
    .B(\soc/cpu/_04679_ ),
    .Y(\soc/cpu/_04680_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09579_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04677_ ),
    .C(\soc/cpu/_04680_ ),
    .Y(\soc/cpu/_00446_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09580_  (.A(\soc/cpu/count_instr[41] ),
    .B(\soc/cpu/_04680_ ),
    .Y(\soc/cpu/_04681_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09581_  (.A(\soc/cpu/count_instr[39] ),
    .B(\soc/cpu/count_instr[40] ),
    .C(net974),
    .D(\soc/cpu/_04675_ ),
    .X(\soc/cpu/_04682_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09582_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04681_ ),
    .C(\soc/cpu/_04682_ ),
    .Y(\soc/cpu/_00447_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09583_  (.A(\soc/cpu/count_instr[34] ),
    .B(\soc/cpu/count_instr[35] ),
    .C(\soc/cpu/count_instr[28] ),
    .X(\soc/cpu/_04683_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09584_  (.A(\soc/cpu/count_instr[32] ),
    .B(\soc/cpu/count_instr[33] ),
    .C(\soc/cpu/count_instr[26] ),
    .D(\soc/cpu/count_instr[27] ),
    .X(\soc/cpu/_04684_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_09585_  (.A(\soc/cpu/count_instr[36] ),
    .B(\soc/cpu/_04662_ ),
    .C(\soc/cpu/_04683_ ),
    .D(\soc/cpu/_04684_ ),
    .Y(\soc/cpu/_04685_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09586_  (.A(\soc/cpu/count_instr[37] ),
    .B(\soc/cpu/count_instr[38] ),
    .Y(\soc/cpu/_04686_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09587_  (.A(\soc/cpu/count_instr[40] ),
    .B(\soc/cpu/count_instr[41] ),
    .Y(\soc/cpu/_04687_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_09588_  (.A(\soc/cpu/_04647_ ),
    .B(\soc/cpu/_04685_ ),
    .C(\soc/cpu/_04686_ ),
    .D(\soc/cpu/_04687_ ),
    .Y(\soc/cpu/_04688_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09589_  (.A(\soc/cpu/count_instr[39] ),
    .B(\soc/cpu/_03995_ ),
    .C(\soc/cpu/_04688_ ),
    .X(\soc/cpu/_04689_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09590_  (.A1(\soc/cpu/count_instr[42] ),
    .A2(\soc/cpu/_04689_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04690_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09591_  (.A1(\soc/cpu/count_instr[42] ),
    .A2(\soc/cpu/_04689_ ),
    .B1(\soc/cpu/_04690_ ),
    .Y(\soc/cpu/_00448_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09592_  (.A1(\soc/cpu/count_instr[42] ),
    .A2(\soc/cpu/_04689_ ),
    .B1(\soc/cpu/count_instr[43] ),
    .Y(\soc/cpu/_04691_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09593_  (.A(net811),
    .B(net792),
    .C(\soc/cpu/_04682_ ),
    .X(\soc/cpu/_04692_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09594_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04691_ ),
    .C(\soc/cpu/_04692_ ),
    .Y(\soc/cpu/_00449_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09595_  (.A1(\soc/cpu/count_instr[44] ),
    .A2(\soc/cpu/_04692_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04693_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09596_  (.A1(\soc/cpu/count_instr[44] ),
    .A2(net812),
    .B1(\soc/cpu/_04693_ ),
    .Y(\soc/cpu/_00450_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09597_  (.A1(\soc/cpu/count_instr[44] ),
    .A2(\soc/cpu/_04692_ ),
    .B1(\soc/cpu/count_instr[45] ),
    .Y(\soc/cpu/_04694_ ));
 sky130_fd_sc_hd__and3_2 \soc/cpu/_09598_  (.A(\soc/cpu/count_instr[44] ),
    .B(\soc/cpu/count_instr[45] ),
    .C(\soc/cpu/_04692_ ),
    .X(\soc/cpu/_04695_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09599_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04694_ ),
    .C(\soc/cpu/_04695_ ),
    .Y(\soc/cpu/_00451_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09600_  (.A1(\soc/cpu/count_instr[46] ),
    .A2(\soc/cpu/_04695_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04696_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09601_  (.A1(\soc/cpu/count_instr[46] ),
    .A2(\soc/cpu/_04695_ ),
    .B1(\soc/cpu/_04696_ ),
    .Y(\soc/cpu/_00452_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09602_  (.A1(\soc/cpu/count_instr[46] ),
    .A2(\soc/cpu/_04695_ ),
    .B1(\soc/cpu/count_instr[47] ),
    .Y(\soc/cpu/_04697_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09603_  (.A(\soc/cpu/count_instr[46] ),
    .B(\soc/cpu/count_instr[47] ),
    .C(\soc/cpu/_04695_ ),
    .X(\soc/cpu/_04698_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09604_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04697_ ),
    .C(\soc/cpu/_04698_ ),
    .Y(\soc/cpu/_00453_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09605_  (.A1(\soc/cpu/count_instr[48] ),
    .A2(\soc/cpu/_04698_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04699_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09606_  (.A(\soc/cpu/count_instr[48] ),
    .B(\soc/cpu/_04698_ ),
    .X(\soc/cpu/_04700_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09607_  (.A(\soc/cpu/_04699_ ),
    .B(\soc/cpu/_04700_ ),
    .Y(\soc/cpu/_00454_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09608_  (.A1(\soc/cpu/count_instr[49] ),
    .A2(\soc/cpu/_04700_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04701_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09609_  (.A(\soc/cpu/count_instr[48] ),
    .B(\soc/cpu/count_instr[49] ),
    .C(\soc/cpu/_04698_ ),
    .X(\soc/cpu/_04702_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09610_  (.A(\soc/cpu/_04701_ ),
    .B(\soc/cpu/_04702_ ),
    .Y(\soc/cpu/_00455_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09611_  (.A1(\soc/cpu/count_instr[50] ),
    .A2(\soc/cpu/_04702_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04703_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09612_  (.A1(\soc/cpu/count_instr[50] ),
    .A2(\soc/cpu/_04702_ ),
    .B1(\soc/cpu/_04703_ ),
    .Y(\soc/cpu/_00456_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09613_  (.A(\soc/cpu/count_instr[50] ),
    .B(\soc/cpu/_04702_ ),
    .Y(\soc/cpu/_04704_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09614_  (.A(\soc/cpu/count_instr[51] ),
    .B(\soc/cpu/_04704_ ),
    .X(\soc/cpu/_04705_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09615_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04705_ ),
    .Y(\soc/cpu/_00457_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09616_  (.A(\soc/cpu/count_instr[41] ),
    .Y(\soc/cpu/_04706_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09617_  (.A(\soc/cpu/count_instr[36] ),
    .B(\soc/cpu/count_instr[37] ),
    .C(\soc/cpu/count_instr[38] ),
    .Y(\soc/cpu/_04707_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09618_  (.A(\soc/cpu/_04706_ ),
    .B(\soc/cpu/_04707_ ),
    .C(\soc/cpu/_04679_ ),
    .Y(\soc/cpu/_04708_ ));
 sky130_fd_sc_hd__nand4_2 \soc/cpu/_09619_  (.A(net811),
    .B(net792),
    .C(\soc/cpu/_04669_ ),
    .D(\soc/cpu/_04708_ ),
    .Y(\soc/cpu/_04709_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09620_  (.A(\soc/cpu/count_instr[47] ),
    .B(\soc/cpu/count_instr[48] ),
    .C(\soc/cpu/count_instr[49] ),
    .Y(\soc/cpu/_04710_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09621_  (.A(\soc/cpu/count_instr[44] ),
    .B(\soc/cpu/count_instr[45] ),
    .C(\soc/cpu/count_instr[50] ),
    .X(\soc/cpu/_04711_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09622_  (.A(\soc/cpu/count_instr[46] ),
    .B(\soc/cpu/count_instr[51] ),
    .C(\soc/cpu/_04711_ ),
    .Y(\soc/cpu/_04712_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09623_  (.A(\soc/cpu/_04709_ ),
    .B(\soc/cpu/_04710_ ),
    .C(\soc/cpu/_04712_ ),
    .Y(\soc/cpu/_04713_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09624_  (.A1(\soc/cpu/count_instr[52] ),
    .A2(\soc/cpu/_04713_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04714_ ));
 sky130_fd_sc_hd__inv_1 \soc/cpu/_09625_  (.A(\soc/cpu/count_instr[52] ),
    .Y(\soc/cpu/_04715_ ));
 sky130_fd_sc_hd__nand3_1 \soc/cpu/_09626_  (.A(\soc/cpu/count_instr[42] ),
    .B(net792),
    .C(\soc/cpu/_04689_ ),
    .Y(\soc/cpu/_04716_ ));
 sky130_fd_sc_hd__nor4_1 \soc/cpu/_09627_  (.A(\soc/cpu/_04715_ ),
    .B(net793),
    .C(\soc/cpu/_04710_ ),
    .D(\soc/cpu/_04712_ ),
    .Y(\soc/cpu/_04717_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09628_  (.A(\soc/cpu/_04714_ ),
    .B(\soc/cpu/_04717_ ),
    .Y(\soc/cpu/_00458_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09629_  (.A1(\soc/cpu/count_instr[53] ),
    .A2(\soc/cpu/_04717_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04718_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09630_  (.A(\soc/cpu/count_instr[52] ),
    .B(\soc/cpu/count_instr[53] ),
    .C(\soc/cpu/_04713_ ),
    .X(\soc/cpu/_04719_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09631_  (.A(\soc/cpu/_04718_ ),
    .B(\soc/cpu/_04719_ ),
    .Y(\soc/cpu/_00459_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09632_  (.A1(\soc/cpu/count_instr[54] ),
    .A2(\soc/cpu/_04719_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04720_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09633_  (.A(\soc/cpu/count_instr[54] ),
    .B(\soc/cpu/_04719_ ),
    .X(\soc/cpu/_04721_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09634_  (.A(\soc/cpu/_04720_ ),
    .B(\soc/cpu/_04721_ ),
    .Y(\soc/cpu/_00460_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09635_  (.A1(\soc/cpu/count_instr[55] ),
    .A2(\soc/cpu/_04721_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04722_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09636_  (.A(\soc/cpu/count_instr[54] ),
    .B(\soc/cpu/count_instr[55] ),
    .C(\soc/cpu/_04719_ ),
    .X(\soc/cpu/_04723_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09637_  (.A(\soc/cpu/_04722_ ),
    .B(\soc/cpu/_04723_ ),
    .Y(\soc/cpu/_00461_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09638_  (.A1(\soc/cpu/count_instr[56] ),
    .A2(\soc/cpu/_04723_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04724_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09639_  (.A(\soc/cpu/count_instr[56] ),
    .B(\soc/cpu/_04723_ ),
    .X(\soc/cpu/_04725_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09640_  (.A(\soc/cpu/_04724_ ),
    .B(\soc/cpu/_04725_ ),
    .Y(\soc/cpu/_00462_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09641_  (.A1(\soc/cpu/count_instr[57] ),
    .A2(\soc/cpu/_04725_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04726_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09642_  (.A(\soc/cpu/count_instr[56] ),
    .B(\soc/cpu/count_instr[57] ),
    .C(\soc/cpu/_04723_ ),
    .X(\soc/cpu/_04727_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09643_  (.A(\soc/cpu/_04726_ ),
    .B(\soc/cpu/_04727_ ),
    .Y(\soc/cpu/_00463_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09644_  (.A1(\soc/cpu/count_instr[58] ),
    .A2(\soc/cpu/_04727_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04728_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09645_  (.A(\soc/cpu/count_instr[46] ),
    .B(\soc/cpu/count_instr[47] ),
    .Y(\soc/cpu/_04729_ ));
 sky130_fd_sc_hd__nand4_1 \soc/cpu/_09646_  (.A(\soc/cpu/count_instr[48] ),
    .B(\soc/cpu/count_instr[49] ),
    .C(\soc/cpu/count_instr[50] ),
    .D(\soc/cpu/count_instr[51] ),
    .Y(\soc/cpu/_04730_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09647_  (.A(\soc/cpu/_04729_ ),
    .B(\soc/cpu/_04730_ ),
    .Y(\soc/cpu/_04731_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09648_  (.A(\soc/cpu/count_instr[52] ),
    .B(\soc/cpu/count_instr[53] ),
    .C(\soc/cpu/_04695_ ),
    .D(\soc/cpu/_04731_ ),
    .X(\soc/cpu/_04732_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09649_  (.A(\soc/cpu/count_instr[54] ),
    .B(\soc/cpu/count_instr[55] ),
    .C(\soc/cpu/_04732_ ),
    .X(\soc/cpu/_04733_ ));
 sky130_fd_sc_hd__and4_1 \soc/cpu/_09650_  (.A(\soc/cpu/count_instr[56] ),
    .B(\soc/cpu/count_instr[57] ),
    .C(\soc/cpu/count_instr[58] ),
    .D(\soc/cpu/_04733_ ),
    .X(\soc/cpu/_04734_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09651_  (.A(\soc/cpu/_04728_ ),
    .B(\soc/cpu/_04734_ ),
    .Y(\soc/cpu/_00464_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09652_  (.A1(\soc/cpu/count_instr[59] ),
    .A2(\soc/cpu/_04734_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04735_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09653_  (.A1(\soc/cpu/count_instr[59] ),
    .A2(\soc/cpu/_04734_ ),
    .B1(\soc/cpu/_04735_ ),
    .Y(\soc/cpu/_00465_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09654_  (.A1(\soc/cpu/count_instr[59] ),
    .A2(\soc/cpu/_04734_ ),
    .B1(\soc/cpu/count_instr[60] ),
    .Y(\soc/cpu/_04736_ ));
 sky130_fd_sc_hd__and3_1 \soc/cpu/_09655_  (.A(\soc/cpu/count_instr[59] ),
    .B(\soc/cpu/count_instr[60] ),
    .C(\soc/cpu/_04734_ ),
    .X(\soc/cpu/_04737_ ));
 sky130_fd_sc_hd__nor3_1 \soc/cpu/_09656_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04736_ ),
    .C(\soc/cpu/_04737_ ),
    .Y(\soc/cpu/_00466_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09657_  (.A1(\soc/cpu/count_instr[61] ),
    .A2(\soc/cpu/_04737_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04738_ ));
 sky130_fd_sc_hd__and2_1 \soc/cpu/_09658_  (.A(\soc/cpu/count_instr[61] ),
    .B(\soc/cpu/_04737_ ),
    .X(\soc/cpu/_04739_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09659_  (.A(\soc/cpu/_04738_ ),
    .B(\soc/cpu/_04739_ ),
    .Y(\soc/cpu/_00467_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09660_  (.A1(\soc/cpu/count_instr[62] ),
    .A2(\soc/cpu/_04739_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04740_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09661_  (.A1(\soc/cpu/count_instr[62] ),
    .A2(\soc/cpu/_04739_ ),
    .B1(\soc/cpu/_04740_ ),
    .Y(\soc/cpu/_00468_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09662_  (.A(\soc/cpu/count_instr[62] ),
    .B(\soc/cpu/_04739_ ),
    .Y(\soc/cpu/_04741_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09663_  (.A(\soc/cpu/count_instr[63] ),
    .B(\soc/cpu/_04741_ ),
    .X(\soc/cpu/_04742_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09664_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04742_ ),
    .Y(\soc/cpu/_00469_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09665_  (.A1(\soc/cpu/irq_state[1] ),
    .A2(\soc/cpu/cpu_state[1] ),
    .B1(\soc/cpu/_03989_ ),
    .Y(\soc/cpu/_04743_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/_09666_  (.A(\soc/cpu/_03397_ ),
    .B(\soc/cpu/_04743_ ),
    .X(\soc/cpu/_04744_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/_09669_  (.A(net413),
    .B(\soc/cpu/_03407_ ),
    .Y(\soc/cpu/_04747_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09671_  (.A1(\soc/cpu/eoi [0]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00785_ ),
    .Y(\soc/cpu/_04749_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09672_  (.A(net131),
    .B(\soc/cpu/_04749_ ),
    .Y(\soc/cpu/_00470_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09674_  (.A1(\soc/cpu/eoi [1]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00753_ ),
    .Y(\soc/cpu/_04751_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09675_  (.A(net132),
    .B(\soc/cpu/_04751_ ),
    .Y(\soc/cpu/_00471_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09676_  (.A1(\soc/cpu/eoi [2]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00762_ ),
    .Y(\soc/cpu/_04752_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09677_  (.A(net132),
    .B(\soc/cpu/_04752_ ),
    .Y(\soc/cpu/_00472_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09678_  (.A1(\soc/cpu/eoi [3]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00771_ ),
    .Y(\soc/cpu/_04753_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09679_  (.A(net131),
    .B(\soc/cpu/_04753_ ),
    .Y(\soc/cpu/_00473_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09680_  (.A1(\soc/cpu/eoi [4]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00759_ ),
    .Y(\soc/cpu/_04754_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09681_  (.A(net131),
    .B(\soc/cpu/_04754_ ),
    .Y(\soc/cpu/_00474_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09682_  (.A1(\soc/cpu/eoi [5]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00754_ ),
    .Y(\soc/cpu/_04755_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09683_  (.A(net132),
    .B(\soc/cpu/_04755_ ),
    .Y(\soc/cpu/_00475_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09684_  (.A1(\soc/cpu/eoi [6]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00776_ ),
    .Y(\soc/cpu/_04756_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09685_  (.A(net132),
    .B(\soc/cpu/_04756_ ),
    .Y(\soc/cpu/_00476_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09686_  (.A1(\soc/cpu/eoi [7]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00758_ ),
    .Y(\soc/cpu/_04757_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09687_  (.A(net131),
    .B(\soc/cpu/_04757_ ),
    .Y(\soc/cpu/_00477_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09688_  (.A1(\soc/cpu/eoi [8]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00765_ ),
    .Y(\soc/cpu/_04758_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09689_  (.A(net131),
    .B(\soc/cpu/_04758_ ),
    .Y(\soc/cpu/_00478_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09690_  (.A1(\soc/cpu/eoi [9]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00774_ ),
    .Y(\soc/cpu/_04759_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09691_  (.A(net131),
    .B(\soc/cpu/_04759_ ),
    .Y(\soc/cpu/_00479_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09694_  (.A1(\soc/cpu/eoi [10]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00748_ ),
    .Y(\soc/cpu/_04762_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09695_  (.A(net131),
    .B(\soc/cpu/_04762_ ),
    .Y(\soc/cpu/_00480_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09697_  (.A1(\soc/cpu/eoi [11]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00784_ ),
    .Y(\soc/cpu/_04764_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09698_  (.A(net131),
    .B(\soc/cpu/_04764_ ),
    .Y(\soc/cpu/_00481_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09699_  (.A1(\soc/cpu/eoi [12]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00755_ ),
    .Y(\soc/cpu/_04765_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09700_  (.A(net131),
    .B(\soc/cpu/_04765_ ),
    .Y(\soc/cpu/_00482_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09701_  (.A1(\soc/cpu/eoi [13]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00786_ ),
    .Y(\soc/cpu/_04766_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09702_  (.A(net131),
    .B(\soc/cpu/_04766_ ),
    .Y(\soc/cpu/_00483_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09703_  (.A1(\soc/cpu/eoi [14]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00763_ ),
    .Y(\soc/cpu/_04767_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09704_  (.A(net131),
    .B(\soc/cpu/_04767_ ),
    .Y(\soc/cpu/_00484_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09705_  (.A1(\soc/cpu/eoi [15]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00773_ ),
    .Y(\soc/cpu/_04768_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09706_  (.A(net131),
    .B(\soc/cpu/_04768_ ),
    .Y(\soc/cpu/_00485_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09707_  (.A1(\soc/cpu/eoi [16]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00781_ ),
    .Y(\soc/cpu/_04769_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09708_  (.A(net131),
    .B(\soc/cpu/_04769_ ),
    .Y(\soc/cpu/_00486_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09709_  (.A1(\soc/cpu/eoi [17]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00770_ ),
    .Y(\soc/cpu/_04770_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09710_  (.A(net131),
    .B(\soc/cpu/_04770_ ),
    .Y(\soc/cpu/_00487_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09711_  (.A1(\soc/cpu/eoi [18]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00750_ ),
    .Y(\soc/cpu/_04771_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09712_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04771_ ),
    .Y(\soc/cpu/_00488_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09713_  (.A1(\soc/cpu/eoi [19]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00779_ ),
    .Y(\soc/cpu/_04772_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09714_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04772_ ),
    .Y(\soc/cpu/_00489_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09717_  (.A1(\soc/cpu/eoi [20]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00749_ ),
    .Y(\soc/cpu/_04775_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09718_  (.A(net131),
    .B(\soc/cpu/_04775_ ),
    .Y(\soc/cpu/_00490_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09720_  (.A1(\soc/cpu/eoi [21]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00764_ ),
    .Y(\soc/cpu/_04777_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09721_  (.A(net131),
    .B(\soc/cpu/_04777_ ),
    .Y(\soc/cpu/_00491_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09722_  (.A1(\soc/cpu/eoi [22]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00783_ ),
    .Y(\soc/cpu/_04778_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09723_  (.A(net131),
    .B(\soc/cpu/_04778_ ),
    .Y(\soc/cpu/_00492_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09724_  (.A1(\soc/cpu/eoi [23]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00768_ ),
    .Y(\soc/cpu/_04779_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09725_  (.A(net131),
    .B(\soc/cpu/_04779_ ),
    .Y(\soc/cpu/_00493_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09726_  (.A1(\soc/cpu/eoi [24]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00780_ ),
    .Y(\soc/cpu/_04780_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09727_  (.A(net131),
    .B(\soc/cpu/_04780_ ),
    .Y(\soc/cpu/_00494_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09728_  (.A1(\soc/cpu/eoi [25]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00752_ ),
    .Y(\soc/cpu/_04781_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09729_  (.A(net131),
    .B(\soc/cpu/_04781_ ),
    .Y(\soc/cpu/_00495_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09730_  (.A1(\soc/cpu/eoi [26]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00775_ ),
    .Y(\soc/cpu/_04782_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09731_  (.A(net131),
    .B(\soc/cpu/_04782_ ),
    .Y(\soc/cpu/_00496_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09732_  (.A1(\soc/cpu/eoi [27]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00760_ ),
    .Y(\soc/cpu/_04783_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09733_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04783_ ),
    .Y(\soc/cpu/_00497_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09734_  (.A1(\soc/cpu/eoi [28]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00757_ ),
    .Y(\soc/cpu/_04784_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09735_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04784_ ),
    .Y(\soc/cpu/_00498_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09736_  (.A1(\soc/cpu/eoi [29]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00747_ ),
    .Y(\soc/cpu/_04785_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09737_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04785_ ),
    .Y(\soc/cpu/_00499_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09738_  (.A1(\soc/cpu/eoi [30]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00769_ ),
    .Y(\soc/cpu/_04786_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09739_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04786_ ),
    .Y(\soc/cpu/_00500_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09741_  (.A1(\soc/cpu/eoi [31]),
    .A2(\soc/cpu/_04744_ ),
    .B1(\soc/cpu/_04747_ ),
    .B2(\soc/cpu/_00778_ ),
    .Y(\soc/cpu/_04788_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09742_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04788_ ),
    .Y(\soc/cpu/_00501_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09743_  (.A(_074_),
    .B(\soc/mem_valid ),
    .Y(\soc/cpu/_04789_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09744_  (.A(\soc/mem_ready ),
    .B(\soc/cpu/_04789_ ),
    .Y(\soc/cpu/_00502_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09745_  (.A(_074_),
    .B(net778),
    .X(\soc/cpu/_00581_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/_09746_  (.A(net413),
    .B(\soc/cpu/instr_timer ),
    .Y(\soc/cpu/_04790_ ));
 sky130_fd_sc_hd__or4_2 \soc/cpu/_09748_  (.A(\soc/cpu/timer[29] ),
    .B(\soc/cpu/timer[28] ),
    .C(\soc/cpu/timer[30] ),
    .D(\soc/cpu/_01014_ ),
    .X(\soc/cpu/_04792_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/cpu/_09749_  (.A1(\soc/cpu/timer[31] ),
    .A2(\soc/cpu/_04792_ ),
    .B1(\soc/cpu/_04790_ ),
    .Y(\soc/cpu/_04793_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09751_  (.A1(\soc/cpu/_02916_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/timer[0] ),
    .X(\soc/cpu/_04795_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09752_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04795_ ),
    .Y(\soc/cpu/_00584_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09753_  (.A(\soc/cpu/timer[1] ),
    .B(net885),
    .X(\soc/cpu/_04796_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09754_  (.A1(\soc/cpu/_02935_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04796_ ),
    .X(\soc/cpu/_04797_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09755_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04797_ ),
    .Y(\soc/cpu/_00585_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09756_  (.A(\soc/cpu/_02945_ ),
    .B(\soc/cpu/_04790_ ),
    .Y(\soc/cpu/_04798_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09757_  (.A1(\soc/cpu/timer[1] ),
    .A2(\soc/cpu/timer[0] ),
    .B1(\soc/cpu/timer[2] ),
    .Y(\soc/cpu/_04799_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09758_  (.A1(\soc/cpu/_00998_ ),
    .A2(\soc/cpu/_04799_ ),
    .B1(\soc/cpu/_04793_ ),
    .Y(\soc/cpu/_04800_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09759_  (.A1(\soc/cpu/_04798_ ),
    .A2(\soc/cpu/_04800_ ),
    .B1(_074_),
    .X(\soc/cpu/_00586_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09760_  (.A(\soc/cpu/timer[3] ),
    .B(\soc/cpu/_00998_ ),
    .X(\soc/cpu/_04801_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09761_  (.A1(\soc/cpu/_02961_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04801_ ),
    .X(\soc/cpu/_04802_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09762_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04802_ ),
    .Y(\soc/cpu/_00587_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09763_  (.A1(\soc/cpu/timer[3] ),
    .A2(\soc/cpu/_00998_ ),
    .B1(\soc/cpu/timer[4] ),
    .X(\soc/cpu/_04803_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09764_  (.A(\soc/cpu/_01028_ ),
    .B(\soc/cpu/_04803_ ),
    .Y(\soc/cpu/_04804_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09765_  (.A1(\soc/cpu/_02980_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04804_ ),
    .X(\soc/cpu/_04805_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09766_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04805_ ),
    .Y(\soc/cpu/_00588_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09767_  (.A1(\soc/cpu/_02987_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01029_ ),
    .X(\soc/cpu/_04806_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09768_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04806_ ),
    .Y(\soc/cpu/_00589_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09769_  (.A1(\soc/cpu/_03008_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01027_ ),
    .X(\soc/cpu/_04807_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09770_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04807_ ),
    .Y(\soc/cpu/_00590_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09771_  (.A(\soc/cpu/timer[7] ),
    .B(\soc/cpu/_01000_ ),
    .Y(\soc/cpu/_04808_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09772_  (.A1(\soc/cpu/_03021_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04808_ ),
    .X(\soc/cpu/_04809_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09773_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04809_ ),
    .Y(\soc/cpu/_00591_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09775_  (.A1(\soc/cpu/_03033_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01026_ ),
    .X(\soc/cpu/_04811_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09776_  (.A(net131),
    .B(\soc/cpu/_04811_ ),
    .Y(\soc/cpu/_00592_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09777_  (.A1(\soc/cpu/_03045_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01025_ ),
    .X(\soc/cpu/_04812_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09778_  (.A(net131),
    .B(\soc/cpu/_04812_ ),
    .Y(\soc/cpu/_00593_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09781_  (.A(\soc/cpu/timer[10] ),
    .B(\soc/cpu/_01002_ ),
    .Y(\soc/cpu/_04815_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09782_  (.A1(\soc/cpu/_03057_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04815_ ),
    .X(\soc/cpu/_04816_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09783_  (.A(net131),
    .B(\soc/cpu/_04816_ ),
    .Y(\soc/cpu/_00594_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09784_  (.A1(\soc/cpu/_03068_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01023_ ),
    .X(\soc/cpu/_04817_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09785_  (.A(net131),
    .B(\soc/cpu/_04817_ ),
    .Y(\soc/cpu/_00595_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09786_  (.A1(\soc/cpu/timer[11] ),
    .A2(\soc/cpu/_01003_ ),
    .B1(\soc/cpu/timer[12] ),
    .X(\soc/cpu/_04818_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09787_  (.A(\soc/cpu/_01004_ ),
    .B(\soc/cpu/_04818_ ),
    .Y(\soc/cpu/_04819_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09788_  (.A1(\soc/cpu/_03076_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04819_ ),
    .X(\soc/cpu/_04820_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09789_  (.A(net131),
    .B(\soc/cpu/_04820_ ),
    .Y(\soc/cpu/_00596_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09790_  (.A(\soc/cpu/timer[13] ),
    .B(\soc/cpu/_01004_ ),
    .Y(\soc/cpu/_04821_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09791_  (.A1(\soc/cpu/_03090_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04821_ ),
    .X(\soc/cpu/_04822_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09792_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04822_ ),
    .Y(\soc/cpu/_00597_ ));
 sky130_fd_sc_hd__nor2b_1 \soc/cpu/_09793_  (.A(\soc/cpu/_01022_ ),
    .B_N(\soc/cpu/_01040_ ),
    .Y(\soc/cpu/_04823_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09794_  (.A1(\soc/cpu/_03102_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04823_ ),
    .X(\soc/cpu/_04824_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09795_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04824_ ),
    .Y(\soc/cpu/_00598_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09796_  (.A(\soc/cpu/timer[15] ),
    .B(\soc/cpu/_01022_ ),
    .Y(\soc/cpu/_04825_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09797_  (.A1(\soc/cpu/_03116_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04825_ ),
    .X(\soc/cpu/_04826_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09798_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04826_ ),
    .Y(\soc/cpu/_00599_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09799_  (.A(\soc/cpu/timer[16] ),
    .B(\soc/cpu/_01006_ ),
    .Y(\soc/cpu/_04827_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09800_  (.A1(\soc/cpu/_03126_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04827_ ),
    .X(\soc/cpu/_04828_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09801_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04828_ ),
    .Y(\soc/cpu/_00600_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09802_  (.A(\soc/cpu/timer[17] ),
    .B(\soc/cpu/_01007_ ),
    .X(\soc/cpu/_04829_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09803_  (.A1(\soc/cpu/_03136_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04829_ ),
    .X(\soc/cpu/_04830_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09804_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04830_ ),
    .Y(\soc/cpu/_00601_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09806_  (.A1(\soc/cpu/timer[17] ),
    .A2(\soc/cpu/_01007_ ),
    .B1(\soc/cpu/timer[18] ),
    .X(\soc/cpu/_04832_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09807_  (.A(\soc/cpu/_01020_ ),
    .B(\soc/cpu/_04832_ ),
    .Y(\soc/cpu/_04833_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09808_  (.A1(\soc/cpu/_03148_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04833_ ),
    .X(\soc/cpu/_04834_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09809_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04834_ ),
    .Y(\soc/cpu/_00602_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09810_  (.A1(\soc/cpu/_03157_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01021_ ),
    .X(\soc/cpu/_04835_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09811_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04835_ ),
    .Y(\soc/cpu/_00603_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09814_  (.A(\soc/cpu/timer[20] ),
    .B(\soc/cpu/_01008_ ),
    .Y(\soc/cpu/_04838_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09815_  (.A1(\soc/cpu/_03170_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04838_ ),
    .X(\soc/cpu/_04839_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09816_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04839_ ),
    .Y(\soc/cpu/_00604_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09817_  (.A(\soc/cpu/_01008_ ),
    .SLEEP(\soc/cpu/timer[20] ),
    .X(\soc/cpu/_04840_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09818_  (.A(\soc/cpu/timer[21] ),
    .B(\soc/cpu/_04840_ ),
    .Y(\soc/cpu/_04841_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09819_  (.A1(\soc/cpu/_03180_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04841_ ),
    .X(\soc/cpu/_04842_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09820_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04842_ ),
    .Y(\soc/cpu/_00605_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09821_  (.A1(\soc/cpu/_03191_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01019_ ),
    .X(\soc/cpu/_04843_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09822_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04843_ ),
    .Y(\soc/cpu/_00606_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/_09823_  (.A1(\soc/cpu/timer[22] ),
    .A2(\soc/cpu/_01010_ ),
    .B1(\soc/cpu/timer[23] ),
    .X(\soc/cpu/_04844_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09824_  (.A(\soc/cpu/_01011_ ),
    .B(\soc/cpu/_04844_ ),
    .Y(\soc/cpu/_04845_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09825_  (.A1(\soc/cpu/_03200_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04845_ ),
    .X(\soc/cpu/_04846_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09826_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04846_ ),
    .Y(\soc/cpu/_00607_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09827_  (.A(\soc/cpu/timer[24] ),
    .B(\soc/cpu/_01011_ ),
    .Y(\soc/cpu/_04847_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09828_  (.A1(\soc/cpu/_03211_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04847_ ),
    .X(\soc/cpu/_04848_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09829_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04848_ ),
    .Y(\soc/cpu/_00608_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09830_  (.A(\soc/cpu/timer[25] ),
    .B(\soc/cpu/_01012_ ),
    .X(\soc/cpu/_04849_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09831_  (.A1(\soc/cpu/_03223_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04849_ ),
    .X(\soc/cpu/_04850_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09832_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04850_ ),
    .Y(\soc/cpu/_00609_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09833_  (.A1(\soc/cpu/_03232_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01018_ ),
    .X(\soc/cpu/_04851_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09834_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04851_ ),
    .Y(\soc/cpu/_00610_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/cpu/_09835_  (.A(\soc/cpu/timer[27] ),
    .B(\soc/cpu/_01013_ ),
    .Y(\soc/cpu/_04852_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09836_  (.A1(\soc/cpu/_03243_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04852_ ),
    .X(\soc/cpu/_04853_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09837_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04853_ ),
    .Y(\soc/cpu/_00611_ ));
 sky130_fd_sc_hd__xor2_1 \soc/cpu/_09838_  (.A(\soc/cpu/timer[28] ),
    .B(\soc/cpu/_01014_ ),
    .X(\soc/cpu/_04854_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09839_  (.A1(\soc/cpu/_03255_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_04854_ ),
    .X(\soc/cpu/_04855_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09840_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04855_ ),
    .Y(\soc/cpu/_00612_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/_09841_  (.A1(\soc/cpu/_03267_ ),
    .A2(\soc/cpu/_04790_ ),
    .B1(\soc/cpu/_04793_ ),
    .B2(\soc/cpu/_01016_ ),
    .X(\soc/cpu/_04856_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09842_  (.A(\soc/cpu/_00840_ ),
    .B(\soc/cpu/_04856_ ),
    .Y(\soc/cpu/_00613_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/_09843_  (.A(\soc/cpu/timer[31] ),
    .SLEEP(\soc/cpu/_04792_ ),
    .X(\soc/cpu/_04857_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/cpu/_09844_  (.A1(\soc/cpu/timer[29] ),
    .A2(\soc/cpu/timer[28] ),
    .A3(\soc/cpu/_01014_ ),
    .B1(\soc/cpu/timer[30] ),
    .Y(\soc/cpu/_04858_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09845_  (.A(\soc/cpu/_04858_ ),
    .B(\soc/cpu/_04790_ ),
    .Y(\soc/cpu/_04859_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09846_  (.A1(\soc/cpu/_04857_ ),
    .A2(\soc/cpu/_04859_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04860_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/cpu/_09847_  (.A1(net414),
    .A2(\soc/cpu/instr_timer ),
    .A3(\soc/cpu/_03277_ ),
    .B1(\soc/cpu/_04860_ ),
    .Y(\soc/cpu/_00614_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/_09848_  (.A(\soc/cpu/timer[31] ),
    .B(\soc/cpu/_04792_ ),
    .Y(\soc/cpu/_04861_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09849_  (.A1(\soc/cpu/cpuregs_rdata1[31] ),
    .A2(\soc/cpu/_02696_ ),
    .B1(\soc/cpu/_04790_ ),
    .Y(\soc/cpu/_04862_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/cpu/_09850_  (.A1(\soc/cpu/_04790_ ),
    .A2(\soc/cpu/_04861_ ),
    .B1(\soc/cpu/_04862_ ),
    .C1(\soc/cpu/_00840_ ),
    .Y(\soc/cpu/_00615_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/_09851_  (.A1(net297),
    .A2(\soc/cpu/_00941_ ),
    .B1(_074_),
    .Y(\soc/cpu/_04863_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09852_  (.A(\soc/cpu/_03370_ ),
    .B(\soc/cpu/_04863_ ),
    .Y(\soc/cpu/_00616_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09853_  (.A1(\soc/cpu/instr_beq ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03353_ ),
    .B2(\soc/cpu/_03365_ ),
    .Y(\soc/cpu/_04864_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09854_  (.A(net132),
    .B(\soc/cpu/_04864_ ),
    .Y(\soc/cpu/_00617_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09855_  (.A1(\soc/cpu/instr_bgeu ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03357_ ),
    .B2(\soc/cpu/_03365_ ),
    .Y(\soc/cpu/_04865_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09856_  (.A(net132),
    .B(\soc/cpu/_04865_ ),
    .Y(\soc/cpu/_00618_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09857_  (.A(\soc/cpu/_02425_ ),
    .B(\soc/cpu/_03341_ ),
    .Y(\soc/cpu/_04866_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/_09858_  (.A1(\soc/cpu/instr_sra ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_04866_ ),
    .Y(\soc/cpu/_04867_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09859_  (.A(net132),
    .B(\soc/cpu/_04867_ ),
    .Y(\soc/cpu/_00621_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/_09860_  (.A1(\soc/cpu/instr_and ),
    .A2(\soc/cpu/_02408_ ),
    .B1(\soc/cpu/_03342_ ),
    .B2(\soc/cpu/_03357_ ),
    .Y(\soc/cpu/_04868_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/_09861_  (.A(net132),
    .B(\soc/cpu/_04868_ ),
    .Y(\soc/cpu/_00622_ ));
 sky130_fd_sc_hd__and2_0 \soc/cpu/_09862_  (.A(_074_),
    .B(\soc/cpu/_00740_ ),
    .X(\soc/cpu/_00665_ ));
 sky130_fd_sc_hd__o211a_1 \soc/cpu/_09863_  (.A1(\soc/cpu/_00839_ ),
    .A2(net154),
    .B1(_074_),
    .C1(\soc/cpu/reg_next_pc[0] ),
    .X(\soc/cpu/_00701_ ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09864_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00064_ ),
    .Q(\soc/cpu/cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09865_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00065_ ),
    .Q(\soc/cpu/cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09866_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00066_ ),
    .Q(\soc/cpu/cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09867_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00067_ ),
    .Q(\soc/cpu/cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09868_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00068_ ),
    .Q(\soc/cpu/cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09869_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00069_ ),
    .Q(\soc/cpu/cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09870_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00070_ ),
    .Q(\soc/cpu/cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09871_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00075_ ),
    .Q(\soc/cpu/mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09872_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00076_ ),
    .Q(\soc/cpu/mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09873_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/cpu/_00077_ ),
    .Q(\soc/cpu/mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09874_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00078_ ),
    .Q(\soc/cpu/mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09875_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/cpu/_00079_ ),
    .Q(\soc/cpu/mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09876_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00080_ ),
    .Q(\soc/cpu/mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09877_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00081_ ),
    .Q(\soc/cpu/mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09878_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00082_ ),
    .Q(\soc/cpu/mem_16bit_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09879_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00083_ ),
    .Q(\soc/cpu/mem_16bit_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09880_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/cpu/_00084_ ),
    .Q(\soc/cpu/mem_16bit_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09881_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00085_ ),
    .Q(\soc/cpu/mem_16bit_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09882_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/cpu/_00086_ ),
    .Q(\soc/cpu/mem_16bit_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09883_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00087_ ),
    .Q(\soc/cpu/mem_16bit_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09884_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00088_ ),
    .Q(\soc/cpu/mem_16bit_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09885_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00089_ ),
    .Q(\soc/cpu/mem_16bit_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09886_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00090_ ),
    .Q(\soc/cpu/mem_16bit_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09887_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00091_ ),
    .Q(\soc/cpu/mem_16bit_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09888_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00092_ ),
    .Q(\soc/cpu/mem_16bit_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09889_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00093_ ),
    .Q(\soc/cpu/mem_16bit_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09890_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00094_ ),
    .Q(\soc/cpu/mem_16bit_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09891_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00095_ ),
    .Q(\soc/cpu/mem_16bit_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09892_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00096_ ),
    .Q(\soc/cpu/mem_16bit_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09893_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00097_ ),
    .Q(\soc/cpu/mem_16bit_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09894_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00058_ ),
    .Q(\soc/cpu/mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09895_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00059_ ),
    .Q(\soc/cpu/mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09896_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00060_ ),
    .Q(\soc/cpu/mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09897_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00036_ ),
    .Q(\soc/cpu/mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09898_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00037_ ),
    .Q(\soc/cpu/mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09899_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00038_ ),
    .Q(\soc/cpu/mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09900_  (.CLK(clknet_leaf_63_clk),
    .D(\soc/cpu/_00039_ ),
    .Q(\soc/cpu/mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09901_  (.CLK(clknet_leaf_63_clk),
    .D(\soc/cpu/_00040_ ),
    .Q(\soc/cpu/mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09902_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00041_ ),
    .Q(\soc/cpu/mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09903_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00042_ ),
    .Q(\soc/cpu/mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09904_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00043_ ),
    .Q(\soc/cpu/mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09905_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00044_ ),
    .Q(\soc/cpu/mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09906_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00045_ ),
    .Q(\soc/cpu/mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09907_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00046_ ),
    .Q(\soc/cpu/mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09908_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00047_ ),
    .Q(\soc/cpu/mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09909_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00048_ ),
    .Q(\soc/cpu/mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09910_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00049_ ),
    .Q(\soc/cpu/mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09911_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00050_ ),
    .Q(\soc/cpu/mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09912_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00051_ ),
    .Q(\soc/cpu/mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09913_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00052_ ),
    .Q(\soc/cpu/mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09914_  (.CLK(clknet_leaf_63_clk),
    .D(\soc/cpu/_00053_ ),
    .Q(\soc/cpu/mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09915_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00054_ ),
    .Q(\soc/cpu/mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09916_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00055_ ),
    .Q(\soc/cpu/mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09917_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00056_ ),
    .Q(\soc/cpu/mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09918_  (.CLK(clknet_leaf_61_clk),
    .D(\soc/cpu/_00057_ ),
    .Q(\soc/cpu/mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09919_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/cpu/_00098_ ),
    .Q(\soc/mem_valid ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09920_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00099_ ),
    .Q(\soc/cpu/prefetched_high_word ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09921_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/cpu/_00100_ ),
    .Q(\soc/cpu/mem_la_secondword ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09922_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00101_ ),
    .Q(\iomem_wstrb[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09923_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00102_ ),
    .Q(\iomem_wstrb[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09924_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00103_ ),
    .Q(\iomem_wstrb[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09925_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00104_ ),
    .Q(\iomem_wstrb[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09926_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00105_ ),
    .Q(\soc/mem_instr ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09927_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00106_ ),
    .Q(\soc/cpu/is_alu_reg_reg ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09928_  (.CLK(clknet_3_3_0_clk),
    .D(\soc/cpu/_00107_ ),
    .Q(\soc/cpu/is_alu_reg_imm ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09929_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00108_ ),
    .Q(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09930_  (.CLK(clknet_leaf_1_clk),
    .D(net752),
    .Q(\soc/cpu/is_sltiu_bltu_sltu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09931_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00034_ ),
    .Q(\soc/cpu/is_slti_blt_slt ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09932_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00109_ ),
    .Q(\soc/cpu/is_slli_srli_srai ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09933_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00110_ ),
    .Q(\soc/cpu/instr_maskirq ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09934_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00111_ ),
    .Q(\soc/cpu/instr_retirq ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09935_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00112_ ),
    .Q(\soc/cpu/decoded_imm_j[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09936_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00113_ ),
    .Q(\soc/cpu/decoded_imm_j[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09937_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00114_ ),
    .Q(\soc/cpu/decoded_imm_j[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09938_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00115_ ),
    .Q(\soc/cpu/decoded_imm_j[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09939_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00116_ ),
    .Q(\soc/cpu/decoded_imm_j[5] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09940_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00117_ ),
    .Q(\soc/cpu/decoded_imm_j[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09941_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00118_ ),
    .Q(\soc/cpu/decoded_imm_j[7] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09942_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00119_ ),
    .Q(\soc/cpu/decoded_imm_j[8] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09943_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00120_ ),
    .Q(\soc/cpu/decoded_imm_j[9] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09944_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00121_ ),
    .Q(\soc/cpu/decoded_imm_j[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09945_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00122_ ),
    .Q(\soc/cpu/decoded_imm_j[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09946_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00123_ ),
    .Q(\soc/cpu/decoded_imm_j[12] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09947_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00124_ ),
    .Q(\soc/cpu/decoded_imm_j[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09948_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00125_ ),
    .Q(\soc/cpu/decoded_imm_j[14] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09949_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00126_ ),
    .Q(\soc/cpu/decoded_imm_j[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09950_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00127_ ),
    .Q(\soc/cpu/decoded_imm_j[16] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09951_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00128_ ),
    .Q(\soc/cpu/decoded_imm_j[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09952_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00129_ ),
    .Q(\soc/cpu/decoded_imm_j[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09953_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00130_ ),
    .Q(\soc/cpu/decoded_imm_j[19] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09954_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00131_ ),
    .Q(\soc/cpu/decoded_imm_j[20] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09955_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00132_ ),
    .Q(\soc/cpu/instr_rdinstrh ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09956_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00133_ ),
    .Q(\soc/cpu/instr_fence ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09957_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00134_ ),
    .Q(\soc/cpu/instr_rdcycleh ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09958_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00135_ ),
    .Q(\soc/cpu/instr_rdcycle ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09959_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00136_ ),
    .Q(\soc/cpu/instr_or ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09960_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00137_ ),
    .Q(\soc/cpu/instr_srl ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09961_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00138_ ),
    .Q(\soc/cpu/instr_xor ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09962_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00139_ ),
    .Q(\soc/cpu/instr_sltu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09963_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00140_ ),
    .Q(\soc/cpu/instr_slt ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09964_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00141_ ),
    .Q(\soc/cpu/instr_sll ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09965_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00142_ ),
    .Q(\soc/cpu/instr_sub ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09966_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00143_ ),
    .Q(\soc/cpu/instr_add ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09967_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00144_ ),
    .Q(\soc/cpu/instr_srli ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09968_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00145_ ),
    .Q(\soc/cpu/instr_slli ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09969_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00146_ ),
    .Q(\soc/cpu/instr_sw ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09970_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00147_ ),
    .Q(\soc/cpu/instr_andi ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09971_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00148_ ),
    .Q(\soc/cpu/instr_ori ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09972_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00149_ ),
    .Q(\soc/cpu/instr_xori ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09973_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00150_ ),
    .Q(\soc/cpu/instr_sltiu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09974_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00151_ ),
    .Q(\soc/cpu/instr_slti ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09975_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00152_ ),
    .Q(\soc/cpu/instr_addi ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09976_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00153_ ),
    .Q(\soc/cpu/instr_sh ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09977_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00154_ ),
    .Q(\soc/cpu/instr_sb ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09978_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00155_ ),
    .Q(\soc/cpu/instr_lhu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09979_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00156_ ),
    .Q(\soc/cpu/instr_lbu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09980_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00157_ ),
    .Q(\soc/cpu/instr_lh ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09981_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00158_ ),
    .Q(\soc/cpu/instr_jalr ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09982_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00159_ ),
    .Q(\soc/cpu/instr_bltu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09983_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00160_ ),
    .Q(\soc/cpu/instr_bge ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09984_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00161_ ),
    .Q(\soc/cpu/instr_blt ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09985_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00162_ ),
    .Q(\soc/cpu/instr_bne ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_09986_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00163_ ),
    .Q(\soc/cpu/instr_jal ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09987_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00164_ ),
    .Q(\soc/cpu/instr_auipc ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09988_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00165_ ),
    .Q(\soc/cpu/do_waitirq ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09989_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/clear_prefetched_high_word ),
    .Q(\soc/cpu/clear_prefetched_high_word_q ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09990_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/alu_out[0] ),
    .Q(\soc/cpu/alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09991_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/alu_out[1] ),
    .Q(\soc/cpu/alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09992_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/alu_out[2] ),
    .Q(\soc/cpu/alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09993_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/alu_out[3] ),
    .Q(\soc/cpu/alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09994_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/alu_out[4] ),
    .Q(\soc/cpu/alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09995_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/alu_out[5] ),
    .Q(\soc/cpu/alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09996_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[6] ),
    .Q(\soc/cpu/alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_09997_  (.CLK(clknet_leaf_94_clk),
    .D(net775),
    .Q(\soc/cpu/alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09998_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[8] ),
    .Q(\soc/cpu/alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_09999_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[9] ),
    .Q(\soc/cpu/alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10000_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[10] ),
    .Q(\soc/cpu/alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10001_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[11] ),
    .Q(\soc/cpu/alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10002_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[12] ),
    .Q(\soc/cpu/alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10003_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/alu_out[13] ),
    .Q(\soc/cpu/alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10004_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/alu_out[14] ),
    .Q(\soc/cpu/alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10005_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/alu_out[15] ),
    .Q(\soc/cpu/alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10006_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/alu_out[16] ),
    .Q(\soc/cpu/alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10007_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/alu_out[17] ),
    .Q(\soc/cpu/alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10008_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/alu_out[18] ),
    .Q(\soc/cpu/alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10009_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[19] ),
    .Q(\soc/cpu/alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10010_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/alu_out[20] ),
    .Q(\soc/cpu/alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10011_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[21] ),
    .Q(\soc/cpu/alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10012_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[22] ),
    .Q(\soc/cpu/alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10013_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[23] ),
    .Q(\soc/cpu/alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10014_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[24] ),
    .Q(\soc/cpu/alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10015_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[25] ),
    .Q(\soc/cpu/alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10016_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[26] ),
    .Q(\soc/cpu/alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10017_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[27] ),
    .Q(\soc/cpu/alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10018_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[28] ),
    .Q(\soc/cpu/alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10019_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[29] ),
    .Q(\soc/cpu/alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10020_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[30] ),
    .Q(\soc/cpu/alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10021_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/alu_out[31] ),
    .Q(\soc/cpu/alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10022_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00166_ ),
    .Q(\soc/cpu/latched_compr ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10023_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00167_ ),
    .Q(\soc/cpu/cpuregs_waddr[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10024_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00168_ ),
    .Q(\soc/cpu/cpuregs_waddr[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10025_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00169_ ),
    .Q(\soc/cpu/cpuregs_waddr[2] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10026_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00170_ ),
    .Q(\soc/cpu/cpuregs_waddr[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10027_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00171_ ),
    .Q(\soc/cpu/cpuregs_waddr[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10028_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00172_ ),
    .Q(\soc/cpu/latched_is_lb ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10029_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00173_ ),
    .Q(\soc/cpu/latched_is_lh ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10030_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00174_ ),
    .Q(\soc/cpu/decoder_pseudo_trigger ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10031_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00175_ ),
    .Q(\soc/cpu/latched_branch ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10032_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00176_ ),
    .Q(\soc/cpu/latched_store ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10033_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00177_ ),
    .Q(\soc/cpu/irq_state[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10034_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00178_ ),
    .Q(\soc/cpu/irq_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10035_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00000_ ),
    .Q(\soc/cpu/decoder_trigger ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10036_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00179_ ),
    .Q(\soc/cpu/mem_do_rinst ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10037_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00180_ ),
    .Q(\soc/cpu/mem_do_prefetch ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10038_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00181_ ),
    .Q(\soc/cpu/reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10039_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00182_ ),
    .Q(\soc/cpu/reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10040_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00183_ ),
    .Q(\soc/cpu/reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10041_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00184_ ),
    .Q(\soc/cpu/reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10042_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00185_ ),
    .Q(\soc/cpu/reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10043_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00186_ ),
    .Q(\soc/cpu/reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10044_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00187_ ),
    .Q(\soc/cpu/reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10045_  (.CLK(clknet_leaf_3_clk),
    .D(net836),
    .Q(\soc/cpu/reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10046_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00189_ ),
    .Q(\soc/cpu/reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10047_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00190_ ),
    .Q(\soc/cpu/reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10048_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00191_ ),
    .Q(\soc/cpu/reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10049_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00192_ ),
    .Q(\soc/cpu/reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10050_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00193_ ),
    .Q(\soc/cpu/reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10051_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00194_ ),
    .Q(\soc/cpu/reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10052_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00195_ ),
    .Q(\soc/cpu/reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10053_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00196_ ),
    .Q(\soc/cpu/reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10054_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00197_ ),
    .Q(\soc/cpu/reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10055_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00198_ ),
    .Q(\soc/cpu/reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10056_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00199_ ),
    .Q(\soc/cpu/reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10057_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00200_ ),
    .Q(\soc/cpu/reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10058_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00201_ ),
    .Q(\soc/cpu/reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10059_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00202_ ),
    .Q(\soc/cpu/reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10060_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00203_ ),
    .Q(\soc/cpu/reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10061_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00204_ ),
    .Q(\soc/cpu/reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10062_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00205_ ),
    .Q(\soc/cpu/reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10063_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00206_ ),
    .Q(\soc/cpu/reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10064_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00207_ ),
    .Q(\soc/cpu/reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10065_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00208_ ),
    .Q(\soc/cpu/reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10066_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00209_ ),
    .Q(\soc/cpu/reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10067_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00210_ ),
    .Q(\soc/cpu/reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10068_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00211_ ),
    .Q(\soc/cpu/reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10069_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00212_ ),
    .Q(\soc/cpu/reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10070_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/_00213_ ),
    .Q(\soc/cpu/irq_mask[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10071_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00214_ ),
    .Q(\soc/cpu/irq_mask[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10072_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00215_ ),
    .Q(\soc/cpu/irq_mask[2] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10073_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00216_ ),
    .Q(\soc/cpu/irq_mask[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10074_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00217_ ),
    .Q(\soc/cpu/irq_mask[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10075_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00218_ ),
    .Q(\soc/cpu/irq_mask[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10076_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00219_ ),
    .Q(\soc/cpu/irq_mask[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10077_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00220_ ),
    .Q(\soc/cpu/irq_mask[7] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10078_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00221_ ),
    .Q(\soc/cpu/irq_mask[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10079_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00222_ ),
    .Q(\soc/cpu/irq_mask[9] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10080_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00223_ ),
    .Q(\soc/cpu/irq_mask[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10081_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00224_ ),
    .Q(\soc/cpu/irq_mask[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10082_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00225_ ),
    .Q(\soc/cpu/irq_mask[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10083_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00226_ ),
    .Q(\soc/cpu/irq_mask[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10084_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00227_ ),
    .Q(\soc/cpu/irq_mask[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10085_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00228_ ),
    .Q(\soc/cpu/irq_mask[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10086_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00229_ ),
    .Q(\soc/cpu/irq_mask[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10087_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00230_ ),
    .Q(\soc/cpu/irq_mask[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10088_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/_00231_ ),
    .Q(\soc/cpu/irq_mask[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10089_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00232_ ),
    .Q(\soc/cpu/irq_mask[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10090_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00233_ ),
    .Q(\soc/cpu/irq_mask[20] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10091_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00234_ ),
    .Q(\soc/cpu/irq_mask[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10092_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00235_ ),
    .Q(\soc/cpu/irq_mask[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10093_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00236_ ),
    .Q(\soc/cpu/irq_mask[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10094_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00237_ ),
    .Q(\soc/cpu/irq_mask[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10095_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00238_ ),
    .Q(\soc/cpu/irq_mask[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10096_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00239_ ),
    .Q(\soc/cpu/irq_mask[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10097_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00240_ ),
    .Q(\soc/cpu/irq_mask[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10098_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00241_ ),
    .Q(\soc/cpu/irq_mask[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10099_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00242_ ),
    .Q(\soc/cpu/irq_mask[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10100_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00243_ ),
    .Q(\soc/cpu/irq_mask[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10101_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00244_ ),
    .Q(\soc/cpu/irq_mask[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10102_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00245_ ),
    .Q(\soc/cpu/irq_active ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10103_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00246_ ),
    .Q(\soc/cpu/irq_delay ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10104_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00247_ ),
    .Q(\soc/cpu/mem_la_wdata [0]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10105_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00248_ ),
    .Q(\soc/cpu/mem_la_wdata [1]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10106_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00249_ ),
    .Q(\soc/cpu/mem_la_wdata [2]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10107_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00250_ ),
    .Q(\soc/cpu/mem_la_wdata [3]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10108_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00251_ ),
    .Q(\soc/cpu/mem_la_wdata [4]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10109_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00252_ ),
    .Q(\soc/cpu/mem_la_wdata [5]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10110_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00253_ ),
    .Q(\soc/cpu/mem_la_wdata [6]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10111_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00254_ ),
    .Q(\soc/cpu/mem_la_wdata [7]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10112_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00255_ ),
    .Q(\soc/cpu/pcpi_rs2 [8]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10113_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00256_ ),
    .Q(\soc/cpu/pcpi_rs2 [9]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10114_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00257_ ),
    .Q(\soc/cpu/pcpi_rs2 [10]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10115_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00258_ ),
    .Q(\soc/cpu/pcpi_rs2 [11]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10116_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00259_ ),
    .Q(\soc/cpu/pcpi_rs2 [12]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10117_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00260_ ),
    .Q(\soc/cpu/pcpi_rs2 [13]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10118_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00261_ ),
    .Q(\soc/cpu/pcpi_rs2 [14]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10119_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00262_ ),
    .Q(\soc/cpu/pcpi_rs2 [15]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10120_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00263_ ),
    .Q(\soc/cpu/pcpi_rs2 [16]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10121_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00264_ ),
    .Q(\soc/cpu/pcpi_rs2 [17]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10122_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00265_ ),
    .Q(\soc/cpu/pcpi_rs2 [18]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10123_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00266_ ),
    .Q(\soc/cpu/pcpi_rs2 [19]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10124_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00267_ ),
    .Q(\soc/cpu/pcpi_rs2 [20]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10125_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00268_ ),
    .Q(\soc/cpu/pcpi_rs2 [21]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10126_  (.CLK(clknet_leaf_11_clk),
    .D(\soc/cpu/_00269_ ),
    .Q(\soc/cpu/pcpi_rs2 [22]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10127_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00270_ ),
    .Q(\soc/cpu/pcpi_rs2 [23]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10128_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00271_ ),
    .Q(\soc/cpu/pcpi_rs2 [24]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10129_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00272_ ),
    .Q(\soc/cpu/pcpi_rs2 [25]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10130_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00273_ ),
    .Q(\soc/cpu/pcpi_rs2 [26]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10131_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00274_ ),
    .Q(\soc/cpu/pcpi_rs2 [27]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10132_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/_00275_ ),
    .Q(\soc/cpu/pcpi_rs2 [28]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10133_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/_00276_ ),
    .Q(\soc/cpu/pcpi_rs2 [29]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10134_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/_00277_ ),
    .Q(\soc/cpu/pcpi_rs2 [30]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10135_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/_00278_ ),
    .Q(\soc/cpu/pcpi_rs2 [31]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10136_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00279_ ),
    .Q(\soc/cpu/pcpi_rs1 [31]));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10137_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00280_ ),
    .Q(\soc/cpu/count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10138_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00281_ ),
    .Q(\soc/cpu/count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10139_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00282_ ),
    .Q(\soc/cpu/count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10140_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00283_ ),
    .Q(\soc/cpu/count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10141_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00284_ ),
    .Q(\soc/cpu/count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10142_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00285_ ),
    .Q(\soc/cpu/count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10143_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00286_ ),
    .Q(\soc/cpu/count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10144_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00287_ ),
    .Q(\soc/cpu/count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10145_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00288_ ),
    .Q(\soc/cpu/count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10146_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00289_ ),
    .Q(\soc/cpu/count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10147_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00290_ ),
    .Q(\soc/cpu/count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10148_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00291_ ),
    .Q(\soc/cpu/count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10149_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00292_ ),
    .Q(\soc/cpu/count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10150_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00293_ ),
    .Q(\soc/cpu/count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10151_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00294_ ),
    .Q(\soc/cpu/count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10152_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00295_ ),
    .Q(\soc/cpu/count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10153_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00296_ ),
    .Q(\soc/cpu/count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10154_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00297_ ),
    .Q(\soc/cpu/count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10155_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00298_ ),
    .Q(\soc/cpu/count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10156_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00299_ ),
    .Q(\soc/cpu/count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10157_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00300_ ),
    .Q(\soc/cpu/count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10158_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00301_ ),
    .Q(\soc/cpu/count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10159_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00302_ ),
    .Q(\soc/cpu/count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10160_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00303_ ),
    .Q(\soc/cpu/count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10161_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00304_ ),
    .Q(\soc/cpu/count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10162_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00305_ ),
    .Q(\soc/cpu/count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10163_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00306_ ),
    .Q(\soc/cpu/count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10164_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00307_ ),
    .Q(\soc/cpu/count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10165_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00308_ ),
    .Q(\soc/cpu/count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10166_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00309_ ),
    .Q(\soc/cpu/count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10167_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00310_ ),
    .Q(\soc/cpu/count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10168_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00311_ ),
    .Q(\soc/cpu/count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10169_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00312_ ),
    .Q(\soc/cpu/count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10170_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00313_ ),
    .Q(\soc/cpu/count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10171_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00314_ ),
    .Q(\soc/cpu/count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10172_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00315_ ),
    .Q(\soc/cpu/count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10173_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00316_ ),
    .Q(\soc/cpu/count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10174_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00317_ ),
    .Q(\soc/cpu/count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10175_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00318_ ),
    .Q(\soc/cpu/count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10176_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00319_ ),
    .Q(\soc/cpu/count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10177_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00320_ ),
    .Q(\soc/cpu/count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10178_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00321_ ),
    .Q(\soc/cpu/count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10179_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00322_ ),
    .Q(\soc/cpu/count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10180_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00323_ ),
    .Q(\soc/cpu/count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10181_  (.CLK(clknet_leaf_54_clk),
    .D(net791),
    .Q(\soc/cpu/count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10182_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00325_ ),
    .Q(\soc/cpu/count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10183_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00326_ ),
    .Q(\soc/cpu/count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10184_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00327_ ),
    .Q(\soc/cpu/count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10185_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00328_ ),
    .Q(\soc/cpu/count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10186_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00329_ ),
    .Q(\soc/cpu/count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10187_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00330_ ),
    .Q(\soc/cpu/count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10188_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00331_ ),
    .Q(\soc/cpu/count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10189_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00332_ ),
    .Q(\soc/cpu/count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10190_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00333_ ),
    .Q(\soc/cpu/count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10191_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00334_ ),
    .Q(\soc/cpu/count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10192_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00335_ ),
    .Q(\soc/cpu/count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10193_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00336_ ),
    .Q(\soc/cpu/count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10194_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00337_ ),
    .Q(\soc/cpu/count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10195_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00338_ ),
    .Q(\soc/cpu/count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10196_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00339_ ),
    .Q(\soc/cpu/count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10197_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00340_ ),
    .Q(\soc/cpu/count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10198_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00341_ ),
    .Q(\soc/cpu/count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10199_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00342_ ),
    .Q(\soc/cpu/count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10200_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00343_ ),
    .Q(\soc/cpu/count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10201_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00344_ ),
    .Q(\soc/cpu/reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10202_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00345_ ),
    .Q(\soc/cpu/reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10203_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00346_ ),
    .Q(\soc/cpu/reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10204_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00347_ ),
    .Q(\soc/cpu/reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10205_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00348_ ),
    .Q(\soc/cpu/reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10206_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00349_ ),
    .Q(\soc/cpu/reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10207_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00350_ ),
    .Q(\soc/cpu/reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10208_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00351_ ),
    .Q(\soc/cpu/reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10209_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00352_ ),
    .Q(\soc/cpu/reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10210_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00353_ ),
    .Q(\soc/cpu/reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10211_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00354_ ),
    .Q(\soc/cpu/reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10212_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00355_ ),
    .Q(\soc/cpu/reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10213_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00356_ ),
    .Q(\soc/cpu/reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10214_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00357_ ),
    .Q(\soc/cpu/reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10215_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00358_ ),
    .Q(\soc/cpu/reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10216_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00359_ ),
    .Q(\soc/cpu/reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10217_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00360_ ),
    .Q(\soc/cpu/reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10218_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00361_ ),
    .Q(\soc/cpu/reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10219_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00362_ ),
    .Q(\soc/cpu/reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10220_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00363_ ),
    .Q(\soc/cpu/reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10221_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00364_ ),
    .Q(\soc/cpu/reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10222_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00365_ ),
    .Q(\soc/cpu/reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10223_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00366_ ),
    .Q(\soc/cpu/reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10224_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00367_ ),
    .Q(\soc/cpu/reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10225_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00368_ ),
    .Q(\soc/cpu/reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10226_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00369_ ),
    .Q(\soc/cpu/reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10227_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00370_ ),
    .Q(\soc/cpu/reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10228_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00371_ ),
    .Q(\soc/cpu/reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10229_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00372_ ),
    .Q(\soc/cpu/reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10230_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00373_ ),
    .Q(\soc/cpu/reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10231_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00374_ ),
    .Q(\soc/cpu/reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10232_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00375_ ),
    .Q(\soc/cpu/reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10233_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00376_ ),
    .Q(\soc/cpu/reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10234_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00377_ ),
    .Q(\soc/cpu/reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10235_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00378_ ),
    .Q(\soc/cpu/reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10236_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00379_ ),
    .Q(\soc/cpu/reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10237_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00380_ ),
    .Q(\soc/cpu/reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10238_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00381_ ),
    .Q(\soc/cpu/reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10239_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00382_ ),
    .Q(\soc/cpu/reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10240_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00383_ ),
    .Q(\soc/cpu/reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10241_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00384_ ),
    .Q(\soc/cpu/reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10242_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00385_ ),
    .Q(\soc/cpu/reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10243_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00386_ ),
    .Q(\soc/cpu/reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10244_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00387_ ),
    .Q(\soc/cpu/reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10245_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00388_ ),
    .Q(\soc/cpu/reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10246_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00389_ ),
    .Q(\soc/cpu/reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10247_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00390_ ),
    .Q(\soc/cpu/reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10248_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00391_ ),
    .Q(\soc/cpu/reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10249_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00392_ ),
    .Q(\soc/cpu/reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10250_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00393_ ),
    .Q(\soc/cpu/reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10251_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00394_ ),
    .Q(\soc/cpu/reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10252_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00395_ ),
    .Q(\soc/cpu/reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10253_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00396_ ),
    .Q(\soc/cpu/reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10254_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00397_ ),
    .Q(\soc/cpu/reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10255_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00398_ ),
    .Q(\soc/cpu/reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10256_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00399_ ),
    .Q(\soc/cpu/reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10257_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00400_ ),
    .Q(\soc/cpu/reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10258_  (.CLK(clknet_leaf_38_clk),
    .D(net820),
    .Q(\soc/cpu/reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10259_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00402_ ),
    .Q(\soc/cpu/reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10260_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00403_ ),
    .Q(\soc/cpu/reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10261_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00404_ ),
    .Q(\soc/cpu/reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10262_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00405_ ),
    .Q(\soc/cpu/reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10263_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00406_ ),
    .Q(\soc/cpu/count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10264_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00407_ ),
    .Q(\soc/cpu/count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10265_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00408_ ),
    .Q(\soc/cpu/count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10266_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00409_ ),
    .Q(\soc/cpu/count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10267_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00410_ ),
    .Q(\soc/cpu/count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10268_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00411_ ),
    .Q(\soc/cpu/count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10269_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00412_ ),
    .Q(\soc/cpu/count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10270_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00413_ ),
    .Q(\soc/cpu/count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10271_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00414_ ),
    .Q(\soc/cpu/count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10272_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00415_ ),
    .Q(\soc/cpu/count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10273_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00416_ ),
    .Q(\soc/cpu/count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10274_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00417_ ),
    .Q(\soc/cpu/count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10275_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00418_ ),
    .Q(\soc/cpu/count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10276_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00419_ ),
    .Q(\soc/cpu/count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10277_  (.CLK(clknet_leaf_54_clk),
    .D(net762),
    .Q(\soc/cpu/count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10278_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00421_ ),
    .Q(\soc/cpu/count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10279_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00422_ ),
    .Q(\soc/cpu/count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10280_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00423_ ),
    .Q(\soc/cpu/count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10281_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00424_ ),
    .Q(\soc/cpu/count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10282_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00425_ ),
    .Q(\soc/cpu/count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10283_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00426_ ),
    .Q(\soc/cpu/count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10284_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00427_ ),
    .Q(\soc/cpu/count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10285_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00428_ ),
    .Q(\soc/cpu/count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10286_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00429_ ),
    .Q(\soc/cpu/count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10287_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00430_ ),
    .Q(\soc/cpu/count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10288_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00431_ ),
    .Q(\soc/cpu/count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10289_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00432_ ),
    .Q(\soc/cpu/count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10290_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00433_ ),
    .Q(\soc/cpu/count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10291_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00434_ ),
    .Q(\soc/cpu/count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10292_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00435_ ),
    .Q(\soc/cpu/count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10293_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00436_ ),
    .Q(\soc/cpu/count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10294_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00437_ ),
    .Q(\soc/cpu/count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10295_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00438_ ),
    .Q(\soc/cpu/count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10296_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00439_ ),
    .Q(\soc/cpu/count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10297_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00440_ ),
    .Q(\soc/cpu/count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10298_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00441_ ),
    .Q(\soc/cpu/count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10299_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00442_ ),
    .Q(\soc/cpu/count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10300_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00443_ ),
    .Q(\soc/cpu/count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10301_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00444_ ),
    .Q(\soc/cpu/count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10302_  (.CLK(clknet_leaf_56_clk),
    .D(\soc/cpu/_00445_ ),
    .Q(\soc/cpu/count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10303_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00446_ ),
    .Q(\soc/cpu/count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10304_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00447_ ),
    .Q(\soc/cpu/count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10305_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00448_ ),
    .Q(\soc/cpu/count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10306_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00449_ ),
    .Q(\soc/cpu/count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10307_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00450_ ),
    .Q(\soc/cpu/count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10308_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00451_ ),
    .Q(\soc/cpu/count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10309_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00452_ ),
    .Q(\soc/cpu/count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10310_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00453_ ),
    .Q(\soc/cpu/count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10311_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00454_ ),
    .Q(\soc/cpu/count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10312_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00455_ ),
    .Q(\soc/cpu/count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10313_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00456_ ),
    .Q(\soc/cpu/count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10314_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00457_ ),
    .Q(\soc/cpu/count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10315_  (.CLK(clknet_leaf_54_clk),
    .D(net794),
    .Q(\soc/cpu/count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10316_  (.CLK(clknet_leaf_54_clk),
    .D(\soc/cpu/_00459_ ),
    .Q(\soc/cpu/count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10317_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00460_ ),
    .Q(\soc/cpu/count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10318_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00461_ ),
    .Q(\soc/cpu/count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10319_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00462_ ),
    .Q(\soc/cpu/count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10320_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00463_ ),
    .Q(\soc/cpu/count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10321_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00464_ ),
    .Q(\soc/cpu/count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10322_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00465_ ),
    .Q(\soc/cpu/count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10323_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00466_ ),
    .Q(\soc/cpu/count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10324_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/_00467_ ),
    .Q(\soc/cpu/count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10325_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00468_ ),
    .Q(\soc/cpu/count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10326_  (.CLK(clknet_leaf_55_clk),
    .D(\soc/cpu/_00469_ ),
    .Q(\soc/cpu/count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10327_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00470_ ),
    .Q(\soc/cpu/eoi [0]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10328_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00471_ ),
    .Q(\soc/cpu/eoi [1]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10329_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00472_ ),
    .Q(\soc/cpu/eoi [2]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10330_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00473_ ),
    .Q(\soc/cpu/eoi [3]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10331_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00474_ ),
    .Q(\soc/cpu/eoi [4]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10332_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00475_ ),
    .Q(\soc/cpu/eoi [5]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10333_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00476_ ),
    .Q(\soc/cpu/eoi [6]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10334_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00477_ ),
    .Q(\soc/cpu/eoi [7]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10335_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00478_ ),
    .Q(\soc/cpu/eoi [8]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10336_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00479_ ),
    .Q(\soc/cpu/eoi [9]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10337_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00480_ ),
    .Q(\soc/cpu/eoi [10]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10338_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00481_ ),
    .Q(\soc/cpu/eoi [11]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10339_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00482_ ),
    .Q(\soc/cpu/eoi [12]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10340_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00483_ ),
    .Q(\soc/cpu/eoi [13]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10341_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00484_ ),
    .Q(\soc/cpu/eoi [14]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10342_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00485_ ),
    .Q(\soc/cpu/eoi [15]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10343_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00486_ ),
    .Q(\soc/cpu/eoi [16]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10344_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00487_ ),
    .Q(\soc/cpu/eoi [17]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10345_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00488_ ),
    .Q(\soc/cpu/eoi [18]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10346_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00489_ ),
    .Q(\soc/cpu/eoi [19]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10347_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00490_ ),
    .Q(\soc/cpu/eoi [20]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10348_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00491_ ),
    .Q(\soc/cpu/eoi [21]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10349_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00492_ ),
    .Q(\soc/cpu/eoi [22]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10350_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00493_ ),
    .Q(\soc/cpu/eoi [23]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10351_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00494_ ),
    .Q(\soc/cpu/eoi [24]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10352_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00495_ ),
    .Q(\soc/cpu/eoi [25]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10353_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00496_ ),
    .Q(\soc/cpu/eoi [26]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10354_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00497_ ),
    .Q(\soc/cpu/eoi [27]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10355_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00498_ ),
    .Q(\soc/cpu/eoi [28]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10356_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00499_ ),
    .Q(\soc/cpu/eoi [29]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10357_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00500_ ),
    .Q(\soc/cpu/eoi [30]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10358_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00501_ ),
    .Q(\soc/cpu/eoi [31]));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10359_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/cpu/_00502_ ),
    .Q(\soc/cpu/last_mem_valid ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10360_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00503_ ),
    .Q(\iomem_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10361_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00504_ ),
    .Q(\iomem_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10362_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00505_ ),
    .Q(\iomem_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10363_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00506_ ),
    .Q(\iomem_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10364_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00507_ ),
    .Q(\iomem_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10365_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00508_ ),
    .Q(\iomem_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10366_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00509_ ),
    .Q(\iomem_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10367_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00510_ ),
    .Q(\iomem_addr[9] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10368_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00511_ ),
    .Q(\iomem_addr[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10369_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00512_ ),
    .Q(\iomem_addr[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10370_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00513_ ),
    .Q(\iomem_addr[12] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10371_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00514_ ),
    .Q(\iomem_addr[13] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10372_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00515_ ),
    .Q(\iomem_addr[14] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10373_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00516_ ),
    .Q(\iomem_addr[15] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10374_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00517_ ),
    .Q(\iomem_addr[16] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10375_  (.CLK(clknet_leaf_90_clk),
    .D(\soc/cpu/_00518_ ),
    .Q(\iomem_addr[17] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10376_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00519_ ),
    .Q(\iomem_addr[18] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10377_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00520_ ),
    .Q(\iomem_addr[19] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10378_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00521_ ),
    .Q(\iomem_addr[20] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10379_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00522_ ),
    .Q(\iomem_addr[21] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10380_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00523_ ),
    .Q(\iomem_addr[22] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10381_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00524_ ),
    .Q(\iomem_addr[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10382_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00525_ ),
    .Q(\iomem_addr[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10383_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00526_ ),
    .Q(\iomem_addr[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10384_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00527_ ),
    .Q(\iomem_addr[26] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10385_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00528_ ),
    .Q(\iomem_addr[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10386_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00529_ ),
    .Q(\iomem_addr[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10387_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00530_ ),
    .Q(\iomem_addr[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10388_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00531_ ),
    .Q(\iomem_addr[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10389_  (.CLK(clknet_leaf_89_clk),
    .D(\soc/cpu/_00532_ ),
    .Q(\iomem_addr[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10390_  (.CLK(clknet_leaf_53_clk),
    .D(\soc/cpu/_00533_ ),
    .Q(\soc/cpu/instr_lui ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10391_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00534_ ),
    .Q(\soc/cpu/instr_srai ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10392_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00535_ ),
    .Q(\soc/cpu/cpuregs_raddr1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10393_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00536_ ),
    .Q(\soc/cpu/cpuregs_raddr1[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10394_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00537_ ),
    .Q(\soc/cpu/cpuregs_raddr1[2] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10395_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00538_ ),
    .Q(\soc/cpu/cpuregs_raddr1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10396_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00539_ ),
    .Q(\soc/cpu/cpuregs_raddr1[4] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10397_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00540_ ),
    .Q(\soc/cpu/cpuregs_raddr2[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10398_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00541_ ),
    .Q(\soc/cpu/cpuregs_raddr2[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10399_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00542_ ),
    .Q(\soc/cpu/cpuregs_raddr2[2] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10400_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00543_ ),
    .Q(\soc/cpu/cpuregs_raddr2[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10401_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00544_ ),
    .Q(\soc/cpu/cpuregs_raddr2[4] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10402_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00545_ ),
    .Q(\soc/cpu/decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10403_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00546_ ),
    .Q(\soc/cpu/decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10404_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00547_ ),
    .Q(\soc/cpu/decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10405_  (.CLK(clknet_leaf_86_clk),
    .D(\soc/cpu/_00548_ ),
    .Q(\soc/cpu/decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10406_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00549_ ),
    .Q(\soc/cpu/decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10407_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00550_ ),
    .Q(\soc/cpu/decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10408_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00551_ ),
    .Q(\soc/cpu/decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10409_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00552_ ),
    .Q(\soc/cpu/decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10410_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00553_ ),
    .Q(\soc/cpu/decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10411_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00554_ ),
    .Q(\soc/cpu/decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10412_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00555_ ),
    .Q(\soc/cpu/decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10413_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00556_ ),
    .Q(\soc/cpu/decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10414_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00557_ ),
    .Q(\soc/cpu/decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10415_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00558_ ),
    .Q(\soc/cpu/decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10416_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00559_ ),
    .Q(\soc/cpu/decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10417_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00560_ ),
    .Q(\soc/cpu/decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10418_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00561_ ),
    .Q(\soc/cpu/decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10419_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00562_ ),
    .Q(\soc/cpu/decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10420_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00563_ ),
    .Q(\soc/cpu/decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10421_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00564_ ),
    .Q(\soc/cpu/decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10422_  (.CLK(clknet_leaf_4_clk),
    .D(\soc/cpu/_00565_ ),
    .Q(\soc/cpu/decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10423_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00566_ ),
    .Q(\soc/cpu/decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10424_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00567_ ),
    .Q(\soc/cpu/decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10425_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00568_ ),
    .Q(\soc/cpu/decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10426_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00569_ ),
    .Q(\soc/cpu/decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10427_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00570_ ),
    .Q(\soc/cpu/decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10428_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00571_ ),
    .Q(\soc/cpu/decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10429_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00572_ ),
    .Q(\soc/cpu/decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10430_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00573_ ),
    .Q(\soc/cpu/decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10431_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00574_ ),
    .Q(\soc/cpu/decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10432_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00575_ ),
    .Q(\soc/cpu/decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10433_  (.CLK(clknet_leaf_40_clk),
    .D(\soc/cpu/_00576_ ),
    .Q(\soc/cpu/decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10434_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00033_ ),
    .Q(\soc/cpu/is_lui_auipc_jal ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10435_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00577_ ),
    .Q(\soc/cpu/is_jalr_addi_slti_sltiu_xori_ori_andi ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10436_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00578_ ),
    .Q(\soc/cpu/is_sb_sh_sw ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10437_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00579_ ),
    .Q(\soc/cpu/is_compare ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10438_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00580_ ),
    .Q(\soc/cpu/compressed_instr ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10439_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00581_ ),
    .Q(\soc/cpu/trap ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10440_  (.CLK(clknet_leaf_38_clk),
    .D(net877),
    .Q(\soc/cpu/irq_pending[0] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10441_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00012_ ),
    .Q(\soc/cpu/irq_pending[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10442_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00023_ ),
    .Q(\soc/cpu/irq_pending[2] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10443_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00026_ ),
    .Q(\soc/cpu/irq_pending[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10444_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00027_ ),
    .Q(\soc/cpu/irq_pending[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10445_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00028_ ),
    .Q(\soc/cpu/irq_pending[5] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10446_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00029_ ),
    .Q(\soc/cpu/irq_pending[6] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10447_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00030_ ),
    .Q(\soc/cpu/irq_pending[7] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10448_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00031_ ),
    .Q(\soc/cpu/irq_pending[8] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10449_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00032_ ),
    .Q(\soc/cpu/irq_pending[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10450_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00002_ ),
    .Q(\soc/cpu/irq_pending[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10451_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00003_ ),
    .Q(\soc/cpu/irq_pending[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10452_  (.CLK(clknet_leaf_5_clk),
    .D(\soc/cpu/_00004_ ),
    .Q(\soc/cpu/irq_pending[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10453_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00005_ ),
    .Q(\soc/cpu/irq_pending[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10454_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00006_ ),
    .Q(\soc/cpu/irq_pending[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10455_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00007_ ),
    .Q(\soc/cpu/irq_pending[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10456_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00008_ ),
    .Q(\soc/cpu/irq_pending[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10457_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00009_ ),
    .Q(\soc/cpu/irq_pending[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10458_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00010_ ),
    .Q(\soc/cpu/irq_pending[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10459_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00011_ ),
    .Q(\soc/cpu/irq_pending[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10460_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00013_ ),
    .Q(\soc/cpu/irq_pending[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10461_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00014_ ),
    .Q(\soc/cpu/irq_pending[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10462_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00015_ ),
    .Q(\soc/cpu/irq_pending[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10463_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00016_ ),
    .Q(\soc/cpu/irq_pending[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10464_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00017_ ),
    .Q(\soc/cpu/irq_pending[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10465_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00018_ ),
    .Q(\soc/cpu/irq_pending[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10466_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00019_ ),
    .Q(\soc/cpu/irq_pending[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10467_  (.CLK(clknet_leaf_39_clk),
    .D(\soc/cpu/_00020_ ),
    .Q(\soc/cpu/irq_pending[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10468_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00021_ ),
    .Q(\soc/cpu/irq_pending[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10469_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00022_ ),
    .Q(\soc/cpu/irq_pending[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10470_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00024_ ),
    .Q(\soc/cpu/irq_pending[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10471_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00025_ ),
    .Q(\soc/cpu/irq_pending[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10472_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00582_ ),
    .Q(\soc/cpu/mem_do_rdata ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10473_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00583_ ),
    .Q(\soc/cpu/mem_do_wdata ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10474_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/_00584_ ),
    .Q(\soc/cpu/timer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10475_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00585_ ),
    .Q(\soc/cpu/timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10476_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00586_ ),
    .Q(\soc/cpu/timer[2] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10477_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00587_ ),
    .Q(\soc/cpu/timer[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10478_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00588_ ),
    .Q(\soc/cpu/timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10479_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00589_ ),
    .Q(\soc/cpu/timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10480_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00590_ ),
    .Q(\soc/cpu/timer[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10481_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/_00591_ ),
    .Q(\soc/cpu/timer[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10482_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00592_ ),
    .Q(\soc/cpu/timer[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10483_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00593_ ),
    .Q(\soc/cpu/timer[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10484_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00594_ ),
    .Q(\soc/cpu/timer[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10485_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00595_ ),
    .Q(\soc/cpu/timer[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10486_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00596_ ),
    .Q(\soc/cpu/timer[12] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10487_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00597_ ),
    .Q(\soc/cpu/timer[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10488_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00598_ ),
    .Q(\soc/cpu/timer[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10489_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00599_ ),
    .Q(\soc/cpu/timer[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10490_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00600_ ),
    .Q(\soc/cpu/timer[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10491_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00601_ ),
    .Q(\soc/cpu/timer[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10492_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/_00602_ ),
    .Q(\soc/cpu/timer[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10493_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00603_ ),
    .Q(\soc/cpu/timer[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10494_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00604_ ),
    .Q(\soc/cpu/timer[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10495_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/_00605_ ),
    .Q(\soc/cpu/timer[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10496_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/_00606_ ),
    .Q(\soc/cpu/timer[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10497_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00607_ ),
    .Q(\soc/cpu/timer[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10498_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00608_ ),
    .Q(\soc/cpu/timer[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10499_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00609_ ),
    .Q(\soc/cpu/timer[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10500_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00610_ ),
    .Q(\soc/cpu/timer[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10501_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/_00611_ ),
    .Q(\soc/cpu/timer[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10502_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/_00612_ ),
    .Q(\soc/cpu/timer[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10503_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/_00613_ ),
    .Q(\soc/cpu/timer[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10504_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00614_ ),
    .Q(\soc/cpu/timer[30] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10505_  (.CLK(clknet_leaf_41_clk),
    .D(\soc/cpu/_00615_ ),
    .Q(\soc/cpu/timer[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10506_  (.CLK(clknet_leaf_59_clk),
    .D(\soc/cpu/_00616_ ),
    .Q(\soc/cpu/latched_stalu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10507_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00617_ ),
    .Q(\soc/cpu/instr_beq ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10508_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00618_ ),
    .Q(\soc/cpu/instr_bgeu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10509_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00619_ ),
    .Q(\soc/cpu/instr_lb ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10510_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00620_ ),
    .Q(\soc/cpu/instr_lw ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10511_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00621_ ),
    .Q(\soc/cpu/instr_sra ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10512_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00622_ ),
    .Q(\soc/cpu/instr_and ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10513_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00623_ ),
    .Q(\soc/cpu/instr_rdinstr ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10514_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00624_ ),
    .Q(\soc/cpu/instr_waitirq ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10515_  (.CLK(clknet_leaf_58_clk),
    .D(\soc/cpu/_00625_ ),
    .Q(\soc/cpu/instr_timer ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10516_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00626_ ),
    .Q(\soc/cpu/decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10517_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00627_ ),
    .Q(\soc/cpu/decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10518_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00628_ ),
    .Q(\soc/cpu/decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10519_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00629_ ),
    .Q(\soc/cpu/decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10520_  (.CLK(clknet_leaf_57_clk),
    .D(\soc/cpu/_00630_ ),
    .Q(\soc/cpu/decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10521_  (.CLK(clknet_leaf_60_clk),
    .D(\soc/cpu/_00631_ ),
    .Q(\soc/cpu/is_lb_lh_lw_lbu_lhu ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10522_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00632_ ),
    .Q(\soc/cpu/is_sll_srl_sra ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10523_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00633_ ),
    .Q(\iomem_wdata[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10524_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00634_ ),
    .Q(\iomem_wdata[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10525_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00635_ ),
    .Q(\iomem_wdata[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10526_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00636_ ),
    .Q(\iomem_wdata[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10527_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00637_ ),
    .Q(\iomem_wdata[4] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10528_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00638_ ),
    .Q(\iomem_wdata[5] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10529_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00639_ ),
    .Q(\iomem_wdata[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10530_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00640_ ),
    .Q(\iomem_wdata[7] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10531_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00641_ ),
    .Q(\iomem_wdata[8] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10532_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00642_ ),
    .Q(\iomem_wdata[9] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10533_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00643_ ),
    .Q(\iomem_wdata[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10534_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00644_ ),
    .Q(\iomem_wdata[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10535_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00645_ ),
    .Q(\iomem_wdata[12] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10536_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00646_ ),
    .Q(\iomem_wdata[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10537_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00647_ ),
    .Q(\iomem_wdata[14] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10538_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00648_ ),
    .Q(\iomem_wdata[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10539_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00649_ ),
    .Q(\iomem_wdata[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10540_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00650_ ),
    .Q(\iomem_wdata[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10541_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00651_ ),
    .Q(\iomem_wdata[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10542_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00652_ ),
    .Q(\iomem_wdata[19] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10543_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00653_ ),
    .Q(\iomem_wdata[20] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10544_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00654_ ),
    .Q(\iomem_wdata[21] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10545_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00655_ ),
    .Q(\iomem_wdata[22] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10546_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00656_ ),
    .Q(\iomem_wdata[23] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10547_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00657_ ),
    .Q(\iomem_wdata[24] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10548_  (.CLK(clknet_leaf_93_clk),
    .D(\soc/cpu/_00658_ ),
    .Q(\iomem_wdata[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10549_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00659_ ),
    .Q(\iomem_wdata[26] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10550_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00660_ ),
    .Q(\iomem_wdata[27] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10551_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00661_ ),
    .Q(\iomem_wdata[28] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10552_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00662_ ),
    .Q(\iomem_wdata[29] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10553_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00663_ ),
    .Q(\iomem_wdata[30] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10554_  (.CLK(clknet_leaf_0_clk),
    .D(\soc/cpu/_00664_ ),
    .Q(\iomem_wdata[31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10555_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/cpu/_00665_ ),
    .Q(\soc/cpu/mem_la_firstword_reg ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10556_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00071_ ),
    .Q(\soc/cpu/mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10557_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00072_ ),
    .Q(\soc/cpu/mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10558_  (.CLK(clknet_leaf_88_clk),
    .D(\soc/cpu/_00073_ ),
    .Q(\soc/cpu/mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10559_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00061_ ),
    .Q(\soc/cpu/reg_sh[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10560_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00062_ ),
    .Q(\soc/cpu/reg_sh[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10561_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00063_ ),
    .Q(\soc/cpu/reg_sh[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10562_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00666_ ),
    .Q(\soc/cpu/mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/cpu/_10563_  (.CLK(clknet_leaf_85_clk),
    .D(\soc/cpu/_00667_ ),
    .Q(\soc/cpu/mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10564_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00668_ ),
    .Q(\soc/cpu/reg_sh[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/_10565_  (.CLK(clknet_leaf_3_clk),
    .D(\soc/cpu/_00669_ ),
    .Q(\soc/cpu/reg_sh[1] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10566_  (.CLK(clknet_leaf_1_clk),
    .D(\soc/cpu/_00670_ ),
    .Q(\soc/cpu/pcpi_rs1 [0]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10567_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00671_ ),
    .Q(\soc/cpu/pcpi_rs1 [1]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10568_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00672_ ),
    .Q(\soc/cpu/pcpi_rs1 [2]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10569_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00673_ ),
    .Q(\soc/cpu/pcpi_rs1 [3]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10570_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00674_ ),
    .Q(\soc/cpu/pcpi_rs1 [4]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10571_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00675_ ),
    .Q(\soc/cpu/pcpi_rs1 [5]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10572_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00676_ ),
    .Q(\soc/cpu/pcpi_rs1 [6]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10573_  (.CLK(clknet_leaf_2_clk),
    .D(\soc/cpu/_00677_ ),
    .Q(\soc/cpu/pcpi_rs1 [7]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10574_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00678_ ),
    .Q(\soc/cpu/pcpi_rs1 [8]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10575_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00679_ ),
    .Q(\soc/cpu/pcpi_rs1 [9]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10576_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00680_ ),
    .Q(\soc/cpu/pcpi_rs1 [10]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10577_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00681_ ),
    .Q(\soc/cpu/pcpi_rs1 [11]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10578_  (.CLK(clknet_leaf_94_clk),
    .D(\soc/cpu/_00682_ ),
    .Q(\soc/cpu/pcpi_rs1 [12]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10579_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00683_ ),
    .Q(\soc/cpu/pcpi_rs1 [13]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10580_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00684_ ),
    .Q(\soc/cpu/pcpi_rs1 [14]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10581_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00685_ ),
    .Q(\soc/cpu/pcpi_rs1 [15]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10582_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00686_ ),
    .Q(\soc/cpu/pcpi_rs1 [16]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10583_  (.CLK(clknet_leaf_10_clk),
    .D(\soc/cpu/_00687_ ),
    .Q(\soc/cpu/pcpi_rs1 [17]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10584_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00688_ ),
    .Q(\soc/cpu/pcpi_rs1 [18]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10585_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00689_ ),
    .Q(\soc/cpu/pcpi_rs1 [19]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10586_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00690_ ),
    .Q(\soc/cpu/pcpi_rs1 [20]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10587_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00691_ ),
    .Q(\soc/cpu/pcpi_rs1 [21]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10588_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00692_ ),
    .Q(\soc/cpu/pcpi_rs1 [22]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10589_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00693_ ),
    .Q(\soc/cpu/pcpi_rs1 [23]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10590_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00694_ ),
    .Q(\soc/cpu/pcpi_rs1 [24]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10591_  (.CLK(clknet_leaf_6_clk),
    .D(\soc/cpu/_00695_ ),
    .Q(\soc/cpu/pcpi_rs1 [25]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10592_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00696_ ),
    .Q(\soc/cpu/pcpi_rs1 [26]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10593_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00697_ ),
    .Q(\soc/cpu/pcpi_rs1 [27]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10594_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00698_ ),
    .Q(\soc/cpu/pcpi_rs1 [28]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10595_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00699_ ),
    .Q(\soc/cpu/pcpi_rs1 [29]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10596_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/_00700_ ),
    .Q(\soc/cpu/pcpi_rs1 [30]));
 sky130_fd_sc_hd__dfxtp_4 \soc/cpu/_10597_  (.CLK(clknet_leaf_87_clk),
    .D(\soc/cpu/_00701_ ),
    .Q(\soc/cpu/reg_next_pc[0] ));
 sky130_fd_sc_hd__conb_1 \soc/_326__458  (.LO(net458));
 sky130_fd_sc_hd__clkinv_16 \soc/cpu/cpuregs/_2520_  (.A(net302),
    .Y(\soc/cpu/cpuregs/_1025_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2530_  (.A0(\soc/cpu/cpuregs/regs[24][0] ),
    .A1(\soc/cpu/cpuregs/regs[25][0] ),
    .A2(\soc/cpu/cpuregs/regs[28][0] ),
    .A3(\soc/cpu/cpuregs/regs[29][0] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1035_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2531_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1035_ ),
    .Y(\soc/cpu/cpuregs/_1036_ ));
 sky130_fd_sc_hd__clkinv_16 \soc/cpu/cpuregs/_2532_  (.A(net313),
    .Y(\soc/cpu/cpuregs/_1037_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2538_  (.A0(\soc/cpu/cpuregs/regs[26][0] ),
    .A1(\soc/cpu/cpuregs/regs[27][0] ),
    .A2(\soc/cpu/cpuregs/regs[30][0] ),
    .A3(\soc/cpu/cpuregs/regs[31][0] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1043_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2541_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1043_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1046_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2548_  (.A0(\soc/cpu/cpuregs/regs[10][0] ),
    .A1(\soc/cpu/cpuregs/regs[11][0] ),
    .A2(\soc/cpu/cpuregs/regs[14][0] ),
    .A3(\soc/cpu/cpuregs/regs[15][0] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1053_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2549_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1053_ ),
    .Y(\soc/cpu/cpuregs/_1054_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2553_  (.A0(\soc/cpu/cpuregs/regs[8][0] ),
    .A1(\soc/cpu/cpuregs/regs[9][0] ),
    .A2(\soc/cpu/cpuregs/regs[12][0] ),
    .A3(\soc/cpu/cpuregs/regs[13][0] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1058_ ));
 sky130_fd_sc_hd__clkinv_16 \soc/cpu/cpuregs/_2554_  (.A(net298),
    .Y(\soc/cpu/cpuregs/_1059_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2556_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1058_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1061_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2557_  (.A1(\soc/cpu/cpuregs/_1036_ ),
    .A2(\soc/cpu/cpuregs/_1046_ ),
    .B1(\soc/cpu/cpuregs/_1054_ ),
    .B2(\soc/cpu/cpuregs/_1061_ ),
    .Y(\soc/cpu/cpuregs/_1062_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2562_  (.A0(\soc/cpu/cpuregs/regs[16][0] ),
    .A1(\soc/cpu/cpuregs/regs[17][0] ),
    .A2(\soc/cpu/cpuregs/regs[20][0] ),
    .A3(\soc/cpu/cpuregs/regs[21][0] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1067_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2563_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1067_ ),
    .Y(\soc/cpu/cpuregs/_1068_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2567_  (.A0(\soc/cpu/cpuregs/regs[18][0] ),
    .A1(\soc/cpu/cpuregs/regs[19][0] ),
    .A2(\soc/cpu/cpuregs/regs[22][0] ),
    .A3(\soc/cpu/cpuregs/regs[23][0] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1072_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2569_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1072_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1074_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2573_  (.A0(\soc/cpu/cpuregs/regs[2][0] ),
    .A1(\soc/cpu/cpuregs/regs[3][0] ),
    .A2(\soc/cpu/cpuregs/regs[6][0] ),
    .A3(\soc/cpu/cpuregs/regs[7][0] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1078_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2574_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1078_ ),
    .Y(\soc/cpu/cpuregs/_1079_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2578_  (.A0(\soc/cpu/cpuregs/regs[0][0] ),
    .A1(\soc/cpu/cpuregs/regs[1][0] ),
    .A2(\soc/cpu/cpuregs/regs[4][0] ),
    .A3(\soc/cpu/cpuregs/regs[5][0] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1083_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2581_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1083_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1086_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2582_  (.A1(\soc/cpu/cpuregs/_1068_ ),
    .A2(\soc/cpu/cpuregs/_1074_ ),
    .B1(\soc/cpu/cpuregs/_1079_ ),
    .B2(\soc/cpu/cpuregs/_1086_ ),
    .C1(\soc/cpu/cpuregs/_1025_ ),
    .Y(\soc/cpu/cpuregs/_1087_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2583_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1062_ ),
    .B1(\soc/cpu/cpuregs/_1087_ ),
    .X(\soc/cpu/cpuregs_rdata2[0] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2585_  (.A0(\soc/cpu/cpuregs/regs[26][1] ),
    .A1(\soc/cpu/cpuregs/regs[27][1] ),
    .A2(\soc/cpu/cpuregs/regs[30][1] ),
    .A3(\soc/cpu/cpuregs/regs[31][1] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1089_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2586_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1089_ ),
    .Y(\soc/cpu/cpuregs/_1090_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2588_  (.A0(\soc/cpu/cpuregs/regs[24][1] ),
    .A1(\soc/cpu/cpuregs/regs[25][1] ),
    .A2(\soc/cpu/cpuregs/regs[28][1] ),
    .A3(\soc/cpu/cpuregs/regs[29][1] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1092_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2589_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1092_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1093_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2592_  (.A0(\soc/cpu/cpuregs/regs[10][1] ),
    .A1(\soc/cpu/cpuregs/regs[11][1] ),
    .A2(\soc/cpu/cpuregs/regs[14][1] ),
    .A3(\soc/cpu/cpuregs/regs[15][1] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1096_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2594_  (.A0(\soc/cpu/cpuregs/regs[8][1] ),
    .A1(\soc/cpu/cpuregs/regs[9][1] ),
    .A2(\soc/cpu/cpuregs/regs[12][1] ),
    .A3(\soc/cpu/cpuregs/regs[13][1] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1098_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2595_  (.A0(\soc/cpu/cpuregs/_1096_ ),
    .A1(\soc/cpu/cpuregs/_1098_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1099_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2597_  (.A1(\soc/cpu/cpuregs/_1090_ ),
    .A2(\soc/cpu/cpuregs/_1093_ ),
    .B1(\soc/cpu/cpuregs/_1099_ ),
    .B2(net300),
    .Y(\soc/cpu/cpuregs/_1101_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2599_  (.A0(\soc/cpu/cpuregs/regs[2][1] ),
    .A1(\soc/cpu/cpuregs/regs[3][1] ),
    .A2(\soc/cpu/cpuregs/regs[6][1] ),
    .A3(\soc/cpu/cpuregs/regs[7][1] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1103_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2600_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1103_ ),
    .Y(\soc/cpu/cpuregs/_1104_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2602_  (.A0(\soc/cpu/cpuregs/regs[0][1] ),
    .A1(\soc/cpu/cpuregs/regs[1][1] ),
    .A2(\soc/cpu/cpuregs/regs[4][1] ),
    .A3(\soc/cpu/cpuregs/regs[5][1] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1106_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2604_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1106_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1108_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2607_  (.A0(\soc/cpu/cpuregs/regs[18][1] ),
    .A1(\soc/cpu/cpuregs/regs[19][1] ),
    .A2(\soc/cpu/cpuregs/regs[22][1] ),
    .A3(\soc/cpu/cpuregs/regs[23][1] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1111_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2610_  (.A0(\soc/cpu/cpuregs/regs[16][1] ),
    .A1(\soc/cpu/cpuregs/regs[17][1] ),
    .A2(\soc/cpu/cpuregs/regs[20][1] ),
    .A3(\soc/cpu/cpuregs/regs[21][1] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1114_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2612_  (.A0(\soc/cpu/cpuregs/_1111_ ),
    .A1(\soc/cpu/cpuregs/_1114_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1116_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2613_  (.A1(\soc/cpu/cpuregs/_1104_ ),
    .A2(\soc/cpu/cpuregs/_1108_ ),
    .B1(\soc/cpu/cpuregs/_1116_ ),
    .B2(\soc/cpu/cpuregs/_1059_ ),
    .C1(\soc/cpu/cpuregs/_1025_ ),
    .Y(\soc/cpu/cpuregs/_1117_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2614_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1101_ ),
    .B1(\soc/cpu/cpuregs/_1117_ ),
    .X(\soc/cpu/cpuregs_rdata2[1] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2616_  (.A0(\soc/cpu/cpuregs/regs[10][2] ),
    .A1(\soc/cpu/cpuregs/regs[11][2] ),
    .A2(\soc/cpu/cpuregs/regs[14][2] ),
    .A3(\soc/cpu/cpuregs/regs[15][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1119_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2617_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1119_ ),
    .Y(\soc/cpu/cpuregs/_1120_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2618_  (.A0(\soc/cpu/cpuregs/regs[8][2] ),
    .A1(\soc/cpu/cpuregs/regs[9][2] ),
    .A2(\soc/cpu/cpuregs/regs[12][2] ),
    .A3(\soc/cpu/cpuregs/regs[13][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1121_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2620_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1121_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1123_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2623_  (.A0(\soc/cpu/cpuregs/regs[24][2] ),
    .A1(\soc/cpu/cpuregs/regs[25][2] ),
    .A2(\soc/cpu/cpuregs/regs[28][2] ),
    .A3(\soc/cpu/cpuregs/regs[29][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1126_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2624_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1126_ ),
    .Y(\soc/cpu/cpuregs/_1127_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2626_  (.A0(\soc/cpu/cpuregs/regs[26][2] ),
    .A1(\soc/cpu/cpuregs/regs[27][2] ),
    .A2(\soc/cpu/cpuregs/regs[30][2] ),
    .A3(\soc/cpu/cpuregs/regs[31][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1129_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2628_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1129_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1131_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2629_  (.A1(\soc/cpu/cpuregs/_1120_ ),
    .A2(\soc/cpu/cpuregs/_1123_ ),
    .B1(\soc/cpu/cpuregs/_1127_ ),
    .B2(\soc/cpu/cpuregs/_1131_ ),
    .Y(\soc/cpu/cpuregs/_1132_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2631_  (.A0(\soc/cpu/cpuregs/regs[2][2] ),
    .A1(\soc/cpu/cpuregs/regs[3][2] ),
    .A2(\soc/cpu/cpuregs/regs[6][2] ),
    .A3(\soc/cpu/cpuregs/regs[7][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1134_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2632_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1134_ ),
    .Y(\soc/cpu/cpuregs/_1135_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2633_  (.A0(\soc/cpu/cpuregs/regs[0][2] ),
    .A1(\soc/cpu/cpuregs/regs[1][2] ),
    .A2(\soc/cpu/cpuregs/regs[4][2] ),
    .A3(\soc/cpu/cpuregs/regs[5][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1136_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2634_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1136_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1137_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2636_  (.A0(\soc/cpu/cpuregs/regs[16][2] ),
    .A1(\soc/cpu/cpuregs/regs[17][2] ),
    .A2(\soc/cpu/cpuregs/regs[20][2] ),
    .A3(\soc/cpu/cpuregs/regs[21][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1139_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2637_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1139_ ),
    .Y(\soc/cpu/cpuregs/_1140_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2639_  (.A0(\soc/cpu/cpuregs/regs[18][2] ),
    .A1(\soc/cpu/cpuregs/regs[19][2] ),
    .A2(\soc/cpu/cpuregs/regs[22][2] ),
    .A3(\soc/cpu/cpuregs/regs[23][2] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1142_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2640_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1142_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1143_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2641_  (.A1(\soc/cpu/cpuregs/_1135_ ),
    .A2(\soc/cpu/cpuregs/_1137_ ),
    .B1(\soc/cpu/cpuregs/_1140_ ),
    .B2(\soc/cpu/cpuregs/_1143_ ),
    .C1(\soc/cpu/cpuregs/_1025_ ),
    .Y(\soc/cpu/cpuregs/_1144_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2642_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1132_ ),
    .B1(\soc/cpu/cpuregs/_1144_ ),
    .X(\soc/cpu/cpuregs_rdata2[2] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2643_  (.A0(\soc/cpu/cpuregs/regs[10][3] ),
    .A1(\soc/cpu/cpuregs/regs[11][3] ),
    .A2(\soc/cpu/cpuregs/regs[14][3] ),
    .A3(\soc/cpu/cpuregs/regs[15][3] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1145_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2644_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1145_ ),
    .Y(\soc/cpu/cpuregs/_1146_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2645_  (.A0(\soc/cpu/cpuregs/regs[8][3] ),
    .A1(\soc/cpu/cpuregs/regs[9][3] ),
    .A2(\soc/cpu/cpuregs/regs[12][3] ),
    .A3(\soc/cpu/cpuregs/regs[13][3] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1147_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2646_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1147_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1148_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2647_  (.A0(\soc/cpu/cpuregs/regs[24][3] ),
    .A1(\soc/cpu/cpuregs/regs[25][3] ),
    .A2(\soc/cpu/cpuregs/regs[28][3] ),
    .A3(\soc/cpu/cpuregs/regs[29][3] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1149_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2648_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1149_ ),
    .Y(\soc/cpu/cpuregs/_1150_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2649_  (.A0(\soc/cpu/cpuregs/regs[26][3] ),
    .A1(\soc/cpu/cpuregs/regs[27][3] ),
    .A2(\soc/cpu/cpuregs/regs[30][3] ),
    .A3(\soc/cpu/cpuregs/regs[31][3] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1151_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2650_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1151_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1152_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2651_  (.A1(\soc/cpu/cpuregs/_1146_ ),
    .A2(\soc/cpu/cpuregs/_1148_ ),
    .B1(\soc/cpu/cpuregs/_1150_ ),
    .B2(\soc/cpu/cpuregs/_1152_ ),
    .Y(\soc/cpu/cpuregs/_1153_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2652_  (.A0(\soc/cpu/cpuregs/regs[2][3] ),
    .A1(\soc/cpu/cpuregs/regs[3][3] ),
    .A2(\soc/cpu/cpuregs/regs[6][3] ),
    .A3(\soc/cpu/cpuregs/regs[7][3] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1154_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2653_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1154_ ),
    .Y(\soc/cpu/cpuregs/_1155_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2654_  (.A0(\soc/cpu/cpuregs/regs[0][3] ),
    .A1(\soc/cpu/cpuregs/regs[1][3] ),
    .A2(\soc/cpu/cpuregs/regs[4][3] ),
    .A3(\soc/cpu/cpuregs/regs[5][3] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1156_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2655_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1156_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1157_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2656_  (.A0(\soc/cpu/cpuregs/regs[16][3] ),
    .A1(\soc/cpu/cpuregs/regs[17][3] ),
    .A2(\soc/cpu/cpuregs/regs[20][3] ),
    .A3(\soc/cpu/cpuregs/regs[21][3] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1158_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2657_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1158_ ),
    .Y(\soc/cpu/cpuregs/_1159_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2658_  (.A0(\soc/cpu/cpuregs/regs[18][3] ),
    .A1(\soc/cpu/cpuregs/regs[19][3] ),
    .A2(\soc/cpu/cpuregs/regs[22][3] ),
    .A3(\soc/cpu/cpuregs/regs[23][3] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1160_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2659_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1160_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1161_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_2660_  (.A1(\soc/cpu/cpuregs/_1155_ ),
    .A2(\soc/cpu/cpuregs/_1157_ ),
    .B1(\soc/cpu/cpuregs/_1159_ ),
    .B2(\soc/cpu/cpuregs/_1161_ ),
    .C1(\soc/cpu/cpuregs/_1025_ ),
    .Y(\soc/cpu/cpuregs/_1162_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2661_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1153_ ),
    .B1(\soc/cpu/cpuregs/_1162_ ),
    .X(\soc/cpu/cpuregs_rdata2[3] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2664_  (.A0(\soc/cpu/cpuregs/regs[26][4] ),
    .A1(\soc/cpu/cpuregs/regs[27][4] ),
    .A2(\soc/cpu/cpuregs/regs[30][4] ),
    .A3(\soc/cpu/cpuregs/regs[31][4] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1165_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2665_  (.A(\soc/cpu/cpuregs/_1025_ ),
    .B(\soc/cpu/cpuregs/_1165_ ),
    .Y(\soc/cpu/cpuregs/_1166_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2667_  (.A0(\soc/cpu/cpuregs/regs[18][4] ),
    .A1(\soc/cpu/cpuregs/regs[19][4] ),
    .A2(\soc/cpu/cpuregs/regs[22][4] ),
    .A3(\soc/cpu/cpuregs/regs[23][4] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1168_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2668_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1168_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1169_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2669_  (.A0(\soc/cpu/cpuregs/regs[2][4] ),
    .A1(\soc/cpu/cpuregs/regs[3][4] ),
    .A2(\soc/cpu/cpuregs/regs[6][4] ),
    .A3(\soc/cpu/cpuregs/regs[7][4] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1170_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2670_  (.A(net303),
    .B(\soc/cpu/cpuregs/_1170_ ),
    .Y(\soc/cpu/cpuregs/_1171_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2671_  (.A0(\soc/cpu/cpuregs/regs[10][4] ),
    .A1(\soc/cpu/cpuregs/regs[11][4] ),
    .A2(\soc/cpu/cpuregs/regs[14][4] ),
    .A3(\soc/cpu/cpuregs/regs[15][4] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1172_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2672_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1172_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1173_ ));
 sky130_fd_sc_hd__o22a_1 \soc/cpu/cpuregs/_2673_  (.A1(\soc/cpu/cpuregs/_1166_ ),
    .A2(\soc/cpu/cpuregs/_1169_ ),
    .B1(\soc/cpu/cpuregs/_1171_ ),
    .B2(\soc/cpu/cpuregs/_1173_ ),
    .X(\soc/cpu/cpuregs/_1174_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2674_  (.A0(\soc/cpu/cpuregs/regs[24][4] ),
    .A1(\soc/cpu/cpuregs/regs[25][4] ),
    .A2(\soc/cpu/cpuregs/regs[28][4] ),
    .A3(\soc/cpu/cpuregs/regs[29][4] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1175_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2676_  (.A0(\soc/cpu/cpuregs/regs[16][4] ),
    .A1(\soc/cpu/cpuregs/regs[17][4] ),
    .A2(\soc/cpu/cpuregs/regs[20][4] ),
    .A3(\soc/cpu/cpuregs/regs[21][4] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1177_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2677_  (.A0(\soc/cpu/cpuregs/regs[8][4] ),
    .A1(\soc/cpu/cpuregs/regs[9][4] ),
    .A2(\soc/cpu/cpuregs/regs[12][4] ),
    .A3(\soc/cpu/cpuregs/regs[13][4] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1178_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2678_  (.A0(\soc/cpu/cpuregs/regs[0][4] ),
    .A1(\soc/cpu/cpuregs/regs[1][4] ),
    .A2(\soc/cpu/cpuregs/regs[4][4] ),
    .A3(\soc/cpu/cpuregs/regs[5][4] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1179_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2679_  (.A0(\soc/cpu/cpuregs/_1175_ ),
    .A1(\soc/cpu/cpuregs/_1177_ ),
    .A2(\soc/cpu/cpuregs/_1178_ ),
    .A3(\soc/cpu/cpuregs/_1179_ ),
    .S0(\soc/cpu/cpuregs/_1025_ ),
    .S1(\soc/cpu/cpuregs/_1059_ ),
    .X(\soc/cpu/cpuregs/_1180_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2680_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1180_ ),
    .Y(\soc/cpu/cpuregs/_1181_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/cpu/cpuregs/_2681_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1174_ ),
    .B1(\soc/cpu/cpuregs/_1181_ ),
    .Y(\soc/cpu/cpuregs_rdata2[4] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2683_  (.A0(\soc/cpu/cpuregs/regs[2][5] ),
    .A1(\soc/cpu/cpuregs/regs[3][5] ),
    .A2(\soc/cpu/cpuregs/regs[6][5] ),
    .A3(\soc/cpu/cpuregs/regs[7][5] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1183_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2684_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1183_ ),
    .Y(\soc/cpu/cpuregs/_1184_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2685_  (.A0(\soc/cpu/cpuregs/regs[0][5] ),
    .A1(\soc/cpu/cpuregs/regs[1][5] ),
    .A2(\soc/cpu/cpuregs/regs[4][5] ),
    .A3(\soc/cpu/cpuregs/regs[5][5] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1185_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2686_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1185_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1186_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2688_  (.A0(\soc/cpu/cpuregs/regs[16][5] ),
    .A1(\soc/cpu/cpuregs/regs[17][5] ),
    .A2(\soc/cpu/cpuregs/regs[20][5] ),
    .A3(\soc/cpu/cpuregs/regs[21][5] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1188_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2689_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1188_ ),
    .Y(\soc/cpu/cpuregs/_1189_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2690_  (.A0(\soc/cpu/cpuregs/regs[18][5] ),
    .A1(\soc/cpu/cpuregs/regs[19][5] ),
    .A2(\soc/cpu/cpuregs/regs[22][5] ),
    .A3(\soc/cpu/cpuregs/regs[23][5] ),
    .S0(net319),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1190_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2691_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1190_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1191_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_2692_  (.A1(\soc/cpu/cpuregs/_1184_ ),
    .A2(\soc/cpu/cpuregs/_1186_ ),
    .B1(\soc/cpu/cpuregs/_1189_ ),
    .B2(\soc/cpu/cpuregs/_1191_ ),
    .Y(\soc/cpu/cpuregs/_1192_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2694_  (.A0(\soc/cpu/cpuregs/regs[10][5] ),
    .A1(\soc/cpu/cpuregs/regs[11][5] ),
    .A2(\soc/cpu/cpuregs/regs[14][5] ),
    .A3(\soc/cpu/cpuregs/regs[15][5] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1194_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2695_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1194_ ),
    .Y(\soc/cpu/cpuregs/_1195_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2696_  (.A0(\soc/cpu/cpuregs/regs[8][5] ),
    .A1(\soc/cpu/cpuregs/regs[9][5] ),
    .A2(\soc/cpu/cpuregs/regs[12][5] ),
    .A3(\soc/cpu/cpuregs/regs[13][5] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1196_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2697_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1196_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1197_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2698_  (.A0(\soc/cpu/cpuregs/regs[24][5] ),
    .A1(\soc/cpu/cpuregs/regs[25][5] ),
    .A2(\soc/cpu/cpuregs/regs[28][5] ),
    .A3(\soc/cpu/cpuregs/regs[29][5] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1198_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2699_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1198_ ),
    .Y(\soc/cpu/cpuregs/_1199_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2700_  (.A0(\soc/cpu/cpuregs/regs[26][5] ),
    .A1(\soc/cpu/cpuregs/regs[27][5] ),
    .A2(\soc/cpu/cpuregs/regs[30][5] ),
    .A3(\soc/cpu/cpuregs/regs[31][5] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1200_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2701_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1200_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1201_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2703_  (.A1(\soc/cpu/cpuregs/_1195_ ),
    .A2(\soc/cpu/cpuregs/_1197_ ),
    .B1(\soc/cpu/cpuregs/_1199_ ),
    .B2(\soc/cpu/cpuregs/_1201_ ),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1203_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2704_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1192_ ),
    .B1(\soc/cpu/cpuregs/_1203_ ),
    .X(\soc/cpu/cpuregs_rdata2[5] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2705_  (.A0(\soc/cpu/cpuregs/regs[16][6] ),
    .A1(\soc/cpu/cpuregs/regs[17][6] ),
    .A2(\soc/cpu/cpuregs/regs[20][6] ),
    .A3(\soc/cpu/cpuregs/regs[21][6] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1204_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2706_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1204_ ),
    .Y(\soc/cpu/cpuregs/_1205_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2708_  (.A0(\soc/cpu/cpuregs/regs[18][6] ),
    .A1(\soc/cpu/cpuregs/regs[19][6] ),
    .A2(\soc/cpu/cpuregs/regs[22][6] ),
    .A3(\soc/cpu/cpuregs/regs[23][6] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1207_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2709_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1207_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1208_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2711_  (.A0(\soc/cpu/cpuregs/regs[2][6] ),
    .A1(\soc/cpu/cpuregs/regs[3][6] ),
    .A2(\soc/cpu/cpuregs/regs[6][6] ),
    .A3(\soc/cpu/cpuregs/regs[7][6] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1210_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2712_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1210_ ),
    .Y(\soc/cpu/cpuregs/_1211_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2714_  (.A0(\soc/cpu/cpuregs/regs[0][6] ),
    .A1(\soc/cpu/cpuregs/regs[1][6] ),
    .A2(\soc/cpu/cpuregs/regs[4][6] ),
    .A3(\soc/cpu/cpuregs/regs[5][6] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1213_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2715_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1213_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1214_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2716_  (.A1(\soc/cpu/cpuregs/_1205_ ),
    .A2(\soc/cpu/cpuregs/_1208_ ),
    .B1(\soc/cpu/cpuregs/_1211_ ),
    .B2(\soc/cpu/cpuregs/_1214_ ),
    .Y(\soc/cpu/cpuregs/_1215_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2717_  (.A0(\soc/cpu/cpuregs/regs[24][6] ),
    .A1(\soc/cpu/cpuregs/regs[25][6] ),
    .A2(\soc/cpu/cpuregs/regs[28][6] ),
    .A3(\soc/cpu/cpuregs/regs[29][6] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1216_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2718_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1216_ ),
    .Y(\soc/cpu/cpuregs/_1217_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2719_  (.A0(\soc/cpu/cpuregs/regs[26][6] ),
    .A1(\soc/cpu/cpuregs/regs[27][6] ),
    .A2(\soc/cpu/cpuregs/regs[30][6] ),
    .A3(\soc/cpu/cpuregs/regs[31][6] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1218_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_2720_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1218_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1219_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2721_  (.A0(\soc/cpu/cpuregs/regs[10][6] ),
    .A1(\soc/cpu/cpuregs/regs[11][6] ),
    .A2(\soc/cpu/cpuregs/regs[14][6] ),
    .A3(\soc/cpu/cpuregs/regs[15][6] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1220_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_2722_  (.A0(\soc/cpu/cpuregs/regs[8][6] ),
    .A1(\soc/cpu/cpuregs/regs[9][6] ),
    .A2(\soc/cpu/cpuregs/regs[12][6] ),
    .A3(\soc/cpu/cpuregs/regs[13][6] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1221_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_2723_  (.A0(\soc/cpu/cpuregs/_1220_ ),
    .A1(\soc/cpu/cpuregs/_1221_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1222_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_2725_  (.A1(\soc/cpu/cpuregs/_1217_ ),
    .A2(\soc/cpu/cpuregs/_1219_ ),
    .B1(\soc/cpu/cpuregs/_1222_ ),
    .B2(net298),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1224_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2726_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1215_ ),
    .B1(\soc/cpu/cpuregs/_1224_ ),
    .X(\soc/cpu/cpuregs_rdata2[6] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2727_  (.A0(\soc/cpu/cpuregs/regs[16][7] ),
    .A1(\soc/cpu/cpuregs/regs[17][7] ),
    .A2(\soc/cpu/cpuregs/regs[20][7] ),
    .A3(\soc/cpu/cpuregs/regs[21][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1225_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2728_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1225_ ),
    .Y(\soc/cpu/cpuregs/_1226_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2729_  (.A0(\soc/cpu/cpuregs/regs[18][7] ),
    .A1(\soc/cpu/cpuregs/regs[19][7] ),
    .A2(\soc/cpu/cpuregs/regs[22][7] ),
    .A3(\soc/cpu/cpuregs/regs[23][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1227_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2730_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1227_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1228_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2731_  (.A0(\soc/cpu/cpuregs/regs[2][7] ),
    .A1(\soc/cpu/cpuregs/regs[3][7] ),
    .A2(\soc/cpu/cpuregs/regs[6][7] ),
    .A3(\soc/cpu/cpuregs/regs[7][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1229_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2732_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1229_ ),
    .Y(\soc/cpu/cpuregs/_1230_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2733_  (.A0(\soc/cpu/cpuregs/regs[0][7] ),
    .A1(\soc/cpu/cpuregs/regs[1][7] ),
    .A2(\soc/cpu/cpuregs/regs[4][7] ),
    .A3(\soc/cpu/cpuregs/regs[5][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1231_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2734_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1231_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1232_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2735_  (.A1(\soc/cpu/cpuregs/_1226_ ),
    .A2(\soc/cpu/cpuregs/_1228_ ),
    .B1(\soc/cpu/cpuregs/_1230_ ),
    .B2(\soc/cpu/cpuregs/_1232_ ),
    .Y(\soc/cpu/cpuregs/_1233_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2736_  (.A0(\soc/cpu/cpuregs/regs[24][7] ),
    .A1(\soc/cpu/cpuregs/regs[25][7] ),
    .A2(\soc/cpu/cpuregs/regs[28][7] ),
    .A3(\soc/cpu/cpuregs/regs[29][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1234_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2737_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1234_ ),
    .Y(\soc/cpu/cpuregs/_1235_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2738_  (.A0(\soc/cpu/cpuregs/regs[26][7] ),
    .A1(\soc/cpu/cpuregs/regs[27][7] ),
    .A2(\soc/cpu/cpuregs/regs[30][7] ),
    .A3(\soc/cpu/cpuregs/regs[31][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1236_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2739_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1236_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1237_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2740_  (.A0(\soc/cpu/cpuregs/regs[10][7] ),
    .A1(\soc/cpu/cpuregs/regs[11][7] ),
    .A2(\soc/cpu/cpuregs/regs[14][7] ),
    .A3(\soc/cpu/cpuregs/regs[15][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1238_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_2741_  (.A0(\soc/cpu/cpuregs/regs[8][7] ),
    .A1(\soc/cpu/cpuregs/regs[9][7] ),
    .A2(\soc/cpu/cpuregs/regs[12][7] ),
    .A3(\soc/cpu/cpuregs/regs[13][7] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1239_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_2742_  (.A0(\soc/cpu/cpuregs/_1238_ ),
    .A1(\soc/cpu/cpuregs/_1239_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1240_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_2743_  (.A1(\soc/cpu/cpuregs/_1235_ ),
    .A2(\soc/cpu/cpuregs/_1237_ ),
    .B1(\soc/cpu/cpuregs/_1240_ ),
    .B2(net298),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1241_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2744_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1233_ ),
    .B1(\soc/cpu/cpuregs/_1241_ ),
    .X(\soc/cpu/cpuregs_rdata2[7] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2746_  (.A0(\soc/cpu/cpuregs/regs[16][8] ),
    .A1(\soc/cpu/cpuregs/regs[17][8] ),
    .A2(\soc/cpu/cpuregs/regs[20][8] ),
    .A3(\soc/cpu/cpuregs/regs[21][8] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1243_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2747_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1243_ ),
    .Y(\soc/cpu/cpuregs/_1244_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2749_  (.A0(\soc/cpu/cpuregs/regs[18][8] ),
    .A1(\soc/cpu/cpuregs/regs[19][8] ),
    .A2(\soc/cpu/cpuregs/regs[22][8] ),
    .A3(\soc/cpu/cpuregs/regs[23][8] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1246_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2750_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1246_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1247_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2751_  (.A0(\soc/cpu/cpuregs/regs[2][8] ),
    .A1(\soc/cpu/cpuregs/regs[3][8] ),
    .A2(\soc/cpu/cpuregs/regs[6][8] ),
    .A3(\soc/cpu/cpuregs/regs[7][8] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1248_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2752_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1248_ ),
    .Y(\soc/cpu/cpuregs/_1249_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2755_  (.A0(\soc/cpu/cpuregs/regs[0][8] ),
    .A1(\soc/cpu/cpuregs/regs[1][8] ),
    .A2(\soc/cpu/cpuregs/regs[4][8] ),
    .A3(\soc/cpu/cpuregs/regs[5][8] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1252_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2756_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1252_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1253_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2757_  (.A1(\soc/cpu/cpuregs/_1244_ ),
    .A2(\soc/cpu/cpuregs/_1247_ ),
    .B1(\soc/cpu/cpuregs/_1249_ ),
    .B2(\soc/cpu/cpuregs/_1253_ ),
    .Y(\soc/cpu/cpuregs/_1254_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2758_  (.A0(\soc/cpu/cpuregs/regs[24][8] ),
    .A1(\soc/cpu/cpuregs/regs[25][8] ),
    .A2(\soc/cpu/cpuregs/regs[28][8] ),
    .A3(\soc/cpu/cpuregs/regs[29][8] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1255_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2759_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1255_ ),
    .Y(\soc/cpu/cpuregs/_1256_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2760_  (.A0(\soc/cpu/cpuregs/regs[26][8] ),
    .A1(\soc/cpu/cpuregs/regs[27][8] ),
    .A2(\soc/cpu/cpuregs/regs[30][8] ),
    .A3(\soc/cpu/cpuregs/regs[31][8] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1257_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2762_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1257_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1259_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2763_  (.A0(\soc/cpu/cpuregs/regs[10][8] ),
    .A1(\soc/cpu/cpuregs/regs[11][8] ),
    .A2(\soc/cpu/cpuregs/regs[14][8] ),
    .A3(\soc/cpu/cpuregs/regs[15][8] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1260_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2764_  (.A0(\soc/cpu/cpuregs/regs[8][8] ),
    .A1(\soc/cpu/cpuregs/regs[9][8] ),
    .A2(\soc/cpu/cpuregs/regs[12][8] ),
    .A3(\soc/cpu/cpuregs/regs[13][8] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1261_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_2765_  (.A0(\soc/cpu/cpuregs/_1260_ ),
    .A1(\soc/cpu/cpuregs/_1261_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1262_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_2766_  (.A1(\soc/cpu/cpuregs/_1256_ ),
    .A2(\soc/cpu/cpuregs/_1259_ ),
    .B1(\soc/cpu/cpuregs/_1262_ ),
    .B2(net298),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1263_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2767_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1254_ ),
    .B1(\soc/cpu/cpuregs/_1263_ ),
    .X(\soc/cpu/cpuregs_rdata2[8] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2770_  (.A0(\soc/cpu/cpuregs/regs[18][9] ),
    .A1(\soc/cpu/cpuregs/regs[19][9] ),
    .A2(\soc/cpu/cpuregs/regs[22][9] ),
    .A3(\soc/cpu/cpuregs/regs[23][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1266_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2772_  (.A0(\soc/cpu/cpuregs/regs[26][9] ),
    .A1(\soc/cpu/cpuregs/regs[27][9] ),
    .A2(\soc/cpu/cpuregs/regs[30][9] ),
    .A3(\soc/cpu/cpuregs/regs[31][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1268_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2773_  (.A0(\soc/cpu/cpuregs/_1266_ ),
    .A1(\soc/cpu/cpuregs/_1268_ ),
    .S(net304),
    .Y(\soc/cpu/cpuregs/_1269_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_2774_  (.A(net301),
    .B(\soc/cpu/cpuregs/_1269_ ),
    .Y(\soc/cpu/cpuregs/_1270_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2775_  (.A0(\soc/cpu/cpuregs/regs[10][9] ),
    .A1(\soc/cpu/cpuregs/regs[11][9] ),
    .A2(\soc/cpu/cpuregs/regs[14][9] ),
    .A3(\soc/cpu/cpuregs/regs[15][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1271_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/cpuregs/_2776_  (.A(\soc/cpu/cpuregs/regs[2][9] ),
    .SLEEP(net308),
    .X(\soc/cpu/cpuregs/_1272_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/cpuregs/_2777_  (.A1(net308),
    .A2(\soc/cpu/cpuregs/regs[6][9] ),
    .B1(\soc/cpu/cpuregs/_1272_ ),
    .C1(net321),
    .X(\soc/cpu/cpuregs/_1273_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2778_  (.A0(\soc/cpu/cpuregs/regs[3][9] ),
    .A1(\soc/cpu/cpuregs/regs[7][9] ),
    .S(net308),
    .Y(\soc/cpu/cpuregs/_1274_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_2779_  (.A1(net321),
    .A2(\soc/cpu/cpuregs/_1274_ ),
    .B1(net304),
    .Y(\soc/cpu/cpuregs/_1275_ ));
 sky130_fd_sc_hd__a221o_1 \soc/cpu/cpuregs/_2781_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1271_ ),
    .B1(\soc/cpu/cpuregs/_1273_ ),
    .B2(\soc/cpu/cpuregs/_1275_ ),
    .C1(net301),
    .X(\soc/cpu/cpuregs/_1277_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2782_  (.A0(\soc/cpu/cpuregs/regs[24][9] ),
    .A1(\soc/cpu/cpuregs/regs[25][9] ),
    .A2(\soc/cpu/cpuregs/regs[28][9] ),
    .A3(\soc/cpu/cpuregs/regs[29][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1278_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2783_  (.A0(\soc/cpu/cpuregs/regs[16][9] ),
    .A1(\soc/cpu/cpuregs/regs[17][9] ),
    .A2(\soc/cpu/cpuregs/regs[20][9] ),
    .A3(\soc/cpu/cpuregs/regs[21][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1279_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2784_  (.A0(\soc/cpu/cpuregs/regs[8][9] ),
    .A1(\soc/cpu/cpuregs/regs[9][9] ),
    .A2(\soc/cpu/cpuregs/regs[12][9] ),
    .A3(\soc/cpu/cpuregs/regs[13][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1280_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2785_  (.A0(\soc/cpu/cpuregs/regs[0][9] ),
    .A1(\soc/cpu/cpuregs/regs[1][9] ),
    .A2(\soc/cpu/cpuregs/regs[4][9] ),
    .A3(\soc/cpu/cpuregs/regs[5][9] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1281_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2786_  (.A0(\soc/cpu/cpuregs/_1278_ ),
    .A1(\soc/cpu/cpuregs/_1279_ ),
    .A2(\soc/cpu/cpuregs/_1280_ ),
    .A3(\soc/cpu/cpuregs/_1281_ ),
    .S0(\soc/cpu/cpuregs/_1025_ ),
    .S1(\soc/cpu/cpuregs/_1059_ ),
    .X(\soc/cpu/cpuregs/_1282_ ));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 \soc/cpu/cpuregs/_2787_  (.A(net153),
    .SLEEP_B(\soc/cpu/cpuregs/_1282_ ),
    .X(\soc/cpu/cpuregs/_1283_ ));
 sky130_fd_sc_hd__a31o_2 \soc/cpu/cpuregs/_2788_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1270_ ),
    .A3(\soc/cpu/cpuregs/_1277_ ),
    .B1(\soc/cpu/cpuregs/_1283_ ),
    .X(\soc/cpu/cpuregs_rdata2[9] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2789_  (.A0(\soc/cpu/cpuregs/regs[2][10] ),
    .A1(\soc/cpu/cpuregs/regs[3][10] ),
    .A2(\soc/cpu/cpuregs/regs[6][10] ),
    .A3(\soc/cpu/cpuregs/regs[7][10] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1284_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2790_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1284_ ),
    .Y(\soc/cpu/cpuregs/_1285_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2791_  (.A0(\soc/cpu/cpuregs/regs[0][10] ),
    .A1(\soc/cpu/cpuregs/regs[1][10] ),
    .A2(\soc/cpu/cpuregs/regs[4][10] ),
    .A3(\soc/cpu/cpuregs/regs[5][10] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1286_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2792_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1286_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1287_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2793_  (.A0(\soc/cpu/cpuregs/regs[16][10] ),
    .A1(\soc/cpu/cpuregs/regs[17][10] ),
    .A2(\soc/cpu/cpuregs/regs[20][10] ),
    .A3(\soc/cpu/cpuregs/regs[21][10] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1288_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2794_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1288_ ),
    .Y(\soc/cpu/cpuregs/_1289_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2795_  (.A0(\soc/cpu/cpuregs/regs[18][10] ),
    .A1(\soc/cpu/cpuregs/regs[19][10] ),
    .A2(\soc/cpu/cpuregs/regs[22][10] ),
    .A3(\soc/cpu/cpuregs/regs[23][10] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1290_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2796_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1290_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1291_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_2797_  (.A1(\soc/cpu/cpuregs/_1285_ ),
    .A2(\soc/cpu/cpuregs/_1287_ ),
    .B1(\soc/cpu/cpuregs/_1289_ ),
    .B2(\soc/cpu/cpuregs/_1291_ ),
    .Y(\soc/cpu/cpuregs/_1292_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2798_  (.A0(\soc/cpu/cpuregs/regs[10][10] ),
    .A1(\soc/cpu/cpuregs/regs[11][10] ),
    .A2(\soc/cpu/cpuregs/regs[14][10] ),
    .A3(\soc/cpu/cpuregs/regs[15][10] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1293_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2799_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1293_ ),
    .Y(\soc/cpu/cpuregs/_1294_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2800_  (.A0(\soc/cpu/cpuregs/regs[8][10] ),
    .A1(\soc/cpu/cpuregs/regs[9][10] ),
    .A2(\soc/cpu/cpuregs/regs[12][10] ),
    .A3(\soc/cpu/cpuregs/regs[13][10] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1295_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2801_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1295_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1296_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2802_  (.A0(\soc/cpu/cpuregs/regs[24][10] ),
    .A1(\soc/cpu/cpuregs/regs[25][10] ),
    .A2(\soc/cpu/cpuregs/regs[28][10] ),
    .A3(\soc/cpu/cpuregs/regs[29][10] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1297_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2803_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1297_ ),
    .Y(\soc/cpu/cpuregs/_1298_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2804_  (.A0(\soc/cpu/cpuregs/regs[26][10] ),
    .A1(\soc/cpu/cpuregs/regs[27][10] ),
    .A2(\soc/cpu/cpuregs/regs[30][10] ),
    .A3(\soc/cpu/cpuregs/regs[31][10] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1299_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2805_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1299_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1300_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2806_  (.A1(\soc/cpu/cpuregs/_1294_ ),
    .A2(\soc/cpu/cpuregs/_1296_ ),
    .B1(\soc/cpu/cpuregs/_1298_ ),
    .B2(\soc/cpu/cpuregs/_1300_ ),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1301_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2807_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1292_ ),
    .B1(\soc/cpu/cpuregs/_1301_ ),
    .X(\soc/cpu/cpuregs_rdata2[10] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2808_  (.A0(\soc/cpu/cpuregs/regs[2][11] ),
    .A1(\soc/cpu/cpuregs/regs[3][11] ),
    .A2(\soc/cpu/cpuregs/regs[6][11] ),
    .A3(\soc/cpu/cpuregs/regs[7][11] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1302_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2810_  (.A0(\soc/cpu/cpuregs/regs[0][11] ),
    .A1(\soc/cpu/cpuregs/regs[1][11] ),
    .A2(\soc/cpu/cpuregs/regs[4][11] ),
    .A3(\soc/cpu/cpuregs/regs[5][11] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1304_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2811_  (.A0(\soc/cpu/cpuregs/_1302_ ),
    .A1(\soc/cpu/cpuregs/_1304_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1305_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2812_  (.A0(\soc/cpu/cpuregs/regs[16][11] ),
    .A1(\soc/cpu/cpuregs/regs[17][11] ),
    .A2(\soc/cpu/cpuregs/regs[20][11] ),
    .A3(\soc/cpu/cpuregs/regs[21][11] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1306_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_2813_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1306_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1307_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2814_  (.A0(\soc/cpu/cpuregs/regs[18][11] ),
    .A1(\soc/cpu/cpuregs/regs[19][11] ),
    .A2(\soc/cpu/cpuregs/regs[22][11] ),
    .A3(\soc/cpu/cpuregs/regs[23][11] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1308_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_2815_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1308_ ),
    .Y(\soc/cpu/cpuregs/_1309_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/cpuregs/_2816_  (.A1(\soc/cpu/cpuregs/_1059_ ),
    .A2(\soc/cpu/cpuregs/_1305_ ),
    .B1(\soc/cpu/cpuregs/_1307_ ),
    .B2(\soc/cpu/cpuregs/_1309_ ),
    .Y(\soc/cpu/cpuregs/_1310_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2818_  (.A0(\soc/cpu/cpuregs/regs[10][11] ),
    .A1(\soc/cpu/cpuregs/regs[11][11] ),
    .A2(\soc/cpu/cpuregs/regs[14][11] ),
    .A3(\soc/cpu/cpuregs/regs[15][11] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1312_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2819_  (.A0(\soc/cpu/cpuregs/regs[8][11] ),
    .A1(\soc/cpu/cpuregs/regs[9][11] ),
    .A2(\soc/cpu/cpuregs/regs[12][11] ),
    .A3(\soc/cpu/cpuregs/regs[13][11] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1313_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2820_  (.A0(\soc/cpu/cpuregs/_1312_ ),
    .A1(\soc/cpu/cpuregs/_1313_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1314_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2821_  (.A0(\soc/cpu/cpuregs/regs[26][11] ),
    .A1(\soc/cpu/cpuregs/regs[27][11] ),
    .A2(\soc/cpu/cpuregs/regs[30][11] ),
    .A3(\soc/cpu/cpuregs/regs[31][11] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1315_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2822_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1315_ ),
    .Y(\soc/cpu/cpuregs/_1316_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2823_  (.A0(\soc/cpu/cpuregs/regs[24][11] ),
    .A1(\soc/cpu/cpuregs/regs[25][11] ),
    .A2(\soc/cpu/cpuregs/regs[28][11] ),
    .A3(\soc/cpu/cpuregs/regs[29][11] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1317_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2824_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1317_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1318_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2825_  (.A1(net299),
    .A2(\soc/cpu/cpuregs/_1314_ ),
    .B1(\soc/cpu/cpuregs/_1316_ ),
    .B2(\soc/cpu/cpuregs/_1318_ ),
    .C1(net302),
    .Y(\soc/cpu/cpuregs/_1319_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2826_  (.A1(net302),
    .A2(\soc/cpu/cpuregs/_1310_ ),
    .B1(\soc/cpu/cpuregs/_1319_ ),
    .X(\soc/cpu/cpuregs_rdata2[11] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2827_  (.A0(\soc/cpu/cpuregs/regs[16][12] ),
    .A1(\soc/cpu/cpuregs/regs[17][12] ),
    .A2(\soc/cpu/cpuregs/regs[20][12] ),
    .A3(\soc/cpu/cpuregs/regs[21][12] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1320_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2828_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1320_ ),
    .Y(\soc/cpu/cpuregs/_1321_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2830_  (.A0(\soc/cpu/cpuregs/regs[18][12] ),
    .A1(\soc/cpu/cpuregs/regs[19][12] ),
    .A2(\soc/cpu/cpuregs/regs[22][12] ),
    .A3(\soc/cpu/cpuregs/regs[23][12] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1323_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2831_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1323_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1324_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2832_  (.A0(\soc/cpu/cpuregs/regs[2][12] ),
    .A1(\soc/cpu/cpuregs/regs[3][12] ),
    .A2(\soc/cpu/cpuregs/regs[6][12] ),
    .A3(\soc/cpu/cpuregs/regs[7][12] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1325_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2833_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1325_ ),
    .Y(\soc/cpu/cpuregs/_1326_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2834_  (.A0(\soc/cpu/cpuregs/regs[0][12] ),
    .A1(\soc/cpu/cpuregs/regs[1][12] ),
    .A2(\soc/cpu/cpuregs/regs[4][12] ),
    .A3(\soc/cpu/cpuregs/regs[5][12] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1327_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2835_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1327_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1328_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2836_  (.A1(\soc/cpu/cpuregs/_1321_ ),
    .A2(\soc/cpu/cpuregs/_1324_ ),
    .B1(\soc/cpu/cpuregs/_1326_ ),
    .B2(\soc/cpu/cpuregs/_1328_ ),
    .Y(\soc/cpu/cpuregs/_1329_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2837_  (.A0(\soc/cpu/cpuregs/regs[24][12] ),
    .A1(\soc/cpu/cpuregs/regs[25][12] ),
    .A2(\soc/cpu/cpuregs/regs[28][12] ),
    .A3(\soc/cpu/cpuregs/regs[29][12] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1330_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2838_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1330_ ),
    .Y(\soc/cpu/cpuregs/_1331_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2839_  (.A0(\soc/cpu/cpuregs/regs[26][12] ),
    .A1(\soc/cpu/cpuregs/regs[27][12] ),
    .A2(\soc/cpu/cpuregs/regs[30][12] ),
    .A3(\soc/cpu/cpuregs/regs[31][12] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1332_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2840_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1332_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1333_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2841_  (.A0(\soc/cpu/cpuregs/regs[10][12] ),
    .A1(\soc/cpu/cpuregs/regs[11][12] ),
    .A2(\soc/cpu/cpuregs/regs[14][12] ),
    .A3(\soc/cpu/cpuregs/regs[15][12] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1334_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2842_  (.A0(\soc/cpu/cpuregs/regs[8][12] ),
    .A1(\soc/cpu/cpuregs/regs[9][12] ),
    .A2(\soc/cpu/cpuregs/regs[12][12] ),
    .A3(\soc/cpu/cpuregs/regs[13][12] ),
    .S0(net321),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1335_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_2844_  (.A0(\soc/cpu/cpuregs/_1334_ ),
    .A1(\soc/cpu/cpuregs/_1335_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1337_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2845_  (.A1(\soc/cpu/cpuregs/_1331_ ),
    .A2(\soc/cpu/cpuregs/_1333_ ),
    .B1(\soc/cpu/cpuregs/_1337_ ),
    .B2(net301),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1338_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_2846_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1329_ ),
    .B1(\soc/cpu/cpuregs/_1338_ ),
    .X(\soc/cpu/cpuregs_rdata2[12] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2848_  (.A0(\soc/cpu/cpuregs/regs[26][13] ),
    .A1(\soc/cpu/cpuregs/regs[27][13] ),
    .A2(\soc/cpu/cpuregs/regs[30][13] ),
    .A3(\soc/cpu/cpuregs/regs[31][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1340_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2849_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1340_ ),
    .Y(\soc/cpu/cpuregs/_1341_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2850_  (.A0(\soc/cpu/cpuregs/regs[24][13] ),
    .A1(\soc/cpu/cpuregs/regs[25][13] ),
    .A2(\soc/cpu/cpuregs/regs[28][13] ),
    .A3(\soc/cpu/cpuregs/regs[29][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1342_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2851_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1342_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1343_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2852_  (.A0(\soc/cpu/cpuregs/regs[10][13] ),
    .A1(\soc/cpu/cpuregs/regs[11][13] ),
    .A2(\soc/cpu/cpuregs/regs[14][13] ),
    .A3(\soc/cpu/cpuregs/regs[15][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1344_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2853_  (.A0(\soc/cpu/cpuregs/regs[8][13] ),
    .A1(\soc/cpu/cpuregs/regs[9][13] ),
    .A2(\soc/cpu/cpuregs/regs[12][13] ),
    .A3(\soc/cpu/cpuregs/regs[13][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1345_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_2854_  (.A0(\soc/cpu/cpuregs/_1344_ ),
    .A1(\soc/cpu/cpuregs/_1345_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1346_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_2855_  (.A1(\soc/cpu/cpuregs/_1341_ ),
    .A2(\soc/cpu/cpuregs/_1343_ ),
    .B1(\soc/cpu/cpuregs/_1346_ ),
    .B2(net298),
    .Y(\soc/cpu/cpuregs/_1347_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2856_  (.A0(\soc/cpu/cpuregs/regs[2][13] ),
    .A1(\soc/cpu/cpuregs/regs[3][13] ),
    .A2(\soc/cpu/cpuregs/regs[6][13] ),
    .A3(\soc/cpu/cpuregs/regs[7][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1348_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2857_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1348_ ),
    .Y(\soc/cpu/cpuregs/_1349_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2860_  (.A0(\soc/cpu/cpuregs/regs[0][13] ),
    .A1(\soc/cpu/cpuregs/regs[1][13] ),
    .A2(\soc/cpu/cpuregs/regs[4][13] ),
    .A3(\soc/cpu/cpuregs/regs[5][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1352_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2861_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1352_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1353_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2862_  (.A0(\soc/cpu/cpuregs/regs[18][13] ),
    .A1(\soc/cpu/cpuregs/regs[19][13] ),
    .A2(\soc/cpu/cpuregs/regs[22][13] ),
    .A3(\soc/cpu/cpuregs/regs[23][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1354_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2863_  (.A0(\soc/cpu/cpuregs/regs[16][13] ),
    .A1(\soc/cpu/cpuregs/regs[17][13] ),
    .A2(\soc/cpu/cpuregs/regs[20][13] ),
    .A3(\soc/cpu/cpuregs/regs[21][13] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1355_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_2864_  (.A0(\soc/cpu/cpuregs/_1354_ ),
    .A1(\soc/cpu/cpuregs/_1355_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1356_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2865_  (.A1(\soc/cpu/cpuregs/_1349_ ),
    .A2(\soc/cpu/cpuregs/_1353_ ),
    .B1(\soc/cpu/cpuregs/_1356_ ),
    .B2(\soc/cpu/cpuregs/_1059_ ),
    .C1(\soc/cpu/cpuregs/_1025_ ),
    .Y(\soc/cpu/cpuregs/_1357_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2866_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1347_ ),
    .B1(\soc/cpu/cpuregs/_1357_ ),
    .X(\soc/cpu/cpuregs_rdata2[13] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2867_  (.A0(\soc/cpu/cpuregs/regs[18][14] ),
    .A1(\soc/cpu/cpuregs/regs[19][14] ),
    .A2(\soc/cpu/cpuregs/regs[22][14] ),
    .A3(\soc/cpu/cpuregs/regs[23][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1358_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2868_  (.A0(\soc/cpu/cpuregs/regs[26][14] ),
    .A1(\soc/cpu/cpuregs/regs[27][14] ),
    .A2(\soc/cpu/cpuregs/regs[30][14] ),
    .A3(\soc/cpu/cpuregs/regs[31][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1359_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2869_  (.A0(\soc/cpu/cpuregs/regs[16][14] ),
    .A1(\soc/cpu/cpuregs/regs[17][14] ),
    .A2(\soc/cpu/cpuregs/regs[20][14] ),
    .A3(\soc/cpu/cpuregs/regs[21][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1360_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2870_  (.A0(\soc/cpu/cpuregs/regs[24][14] ),
    .A1(\soc/cpu/cpuregs/regs[25][14] ),
    .A2(\soc/cpu/cpuregs/regs[28][14] ),
    .A3(\soc/cpu/cpuregs/regs[29][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1361_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2871_  (.A0(\soc/cpu/cpuregs/_1358_ ),
    .A1(\soc/cpu/cpuregs/_1359_ ),
    .A2(\soc/cpu/cpuregs/_1360_ ),
    .A3(\soc/cpu/cpuregs/_1361_ ),
    .S0(net302),
    .S1(\soc/cpu/cpuregs/_1037_ ),
    .X(\soc/cpu/cpuregs/_1362_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_2872_  (.A(\soc/cpu/cpuregs/_1059_ ),
    .B(\soc/cpu/cpuregs/_1362_ ),
    .Y(\soc/cpu/cpuregs/_1363_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2873_  (.A0(\soc/cpu/cpuregs/regs[2][14] ),
    .A1(\soc/cpu/cpuregs/regs[3][14] ),
    .A2(\soc/cpu/cpuregs/regs[6][14] ),
    .A3(\soc/cpu/cpuregs/regs[7][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1364_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2874_  (.A0(\soc/cpu/cpuregs/regs[10][14] ),
    .A1(\soc/cpu/cpuregs/regs[11][14] ),
    .A2(\soc/cpu/cpuregs/regs[14][14] ),
    .A3(\soc/cpu/cpuregs/regs[15][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1365_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2875_  (.A0(\soc/cpu/cpuregs/regs[0][14] ),
    .A1(\soc/cpu/cpuregs/regs[1][14] ),
    .A2(\soc/cpu/cpuregs/regs[4][14] ),
    .A3(\soc/cpu/cpuregs/regs[5][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1366_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2876_  (.A0(\soc/cpu/cpuregs/regs[8][14] ),
    .A1(\soc/cpu/cpuregs/regs[9][14] ),
    .A2(\soc/cpu/cpuregs/regs[12][14] ),
    .A3(\soc/cpu/cpuregs/regs[13][14] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1367_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2877_  (.A0(\soc/cpu/cpuregs/_1364_ ),
    .A1(\soc/cpu/cpuregs/_1365_ ),
    .A2(\soc/cpu/cpuregs/_1366_ ),
    .A3(\soc/cpu/cpuregs/_1367_ ),
    .S0(net302),
    .S1(\soc/cpu/cpuregs/_1037_ ),
    .X(\soc/cpu/cpuregs/_1368_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_2878_  (.A(net300),
    .B(\soc/cpu/cpuregs/_1368_ ),
    .Y(\soc/cpu/cpuregs/_1369_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_2879_  (.A(\soc/cpu/cpuregs/_1363_ ),
    .B(\soc/cpu/cpuregs/_1369_ ),
    .Y(\soc/cpu/cpuregs_rdata2[14] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2880_  (.A0(\soc/cpu/cpuregs/regs[10][15] ),
    .A1(\soc/cpu/cpuregs/regs[11][15] ),
    .A2(\soc/cpu/cpuregs/regs[14][15] ),
    .A3(\soc/cpu/cpuregs/regs[15][15] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1370_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2881_  (.A0(\soc/cpu/cpuregs/regs[2][15] ),
    .A1(\soc/cpu/cpuregs/regs[3][15] ),
    .A2(\soc/cpu/cpuregs/regs[6][15] ),
    .A3(\soc/cpu/cpuregs/regs[7][15] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1371_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2882_  (.A0(\soc/cpu/cpuregs/regs[26][15] ),
    .A1(\soc/cpu/cpuregs/regs[27][15] ),
    .A2(\soc/cpu/cpuregs/regs[30][15] ),
    .A3(\soc/cpu/cpuregs/regs[31][15] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1372_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2883_  (.A0(\soc/cpu/cpuregs/regs[18][15] ),
    .A1(\soc/cpu/cpuregs/regs[19][15] ),
    .A2(\soc/cpu/cpuregs/regs[22][15] ),
    .A3(\soc/cpu/cpuregs/regs[23][15] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1373_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2884_  (.A0(\soc/cpu/cpuregs/_1370_ ),
    .A1(\soc/cpu/cpuregs/_1371_ ),
    .A2(\soc/cpu/cpuregs/_1372_ ),
    .A3(\soc/cpu/cpuregs/_1373_ ),
    .S0(\soc/cpu/cpuregs/_1025_ ),
    .S1(net298),
    .X(\soc/cpu/cpuregs/_1374_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2885_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1374_ ),
    .Y(\soc/cpu/cpuregs/_1375_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2886_  (.A0(\soc/cpu/cpuregs/regs[24][15] ),
    .A1(\soc/cpu/cpuregs/regs[25][15] ),
    .A2(\soc/cpu/cpuregs/regs[28][15] ),
    .A3(\soc/cpu/cpuregs/regs[29][15] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1376_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2887_  (.A0(\soc/cpu/cpuregs/regs[16][15] ),
    .A1(\soc/cpu/cpuregs/regs[17][15] ),
    .A2(\soc/cpu/cpuregs/regs[20][15] ),
    .A3(\soc/cpu/cpuregs/regs[21][15] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1377_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2888_  (.A0(\soc/cpu/cpuregs/regs[8][15] ),
    .A1(\soc/cpu/cpuregs/regs[9][15] ),
    .A2(\soc/cpu/cpuregs/regs[12][15] ),
    .A3(\soc/cpu/cpuregs/regs[13][15] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1378_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2889_  (.A0(\soc/cpu/cpuregs/regs[0][15] ),
    .A1(\soc/cpu/cpuregs/regs[1][15] ),
    .A2(\soc/cpu/cpuregs/regs[4][15] ),
    .A3(\soc/cpu/cpuregs/regs[5][15] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1379_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2890_  (.A0(\soc/cpu/cpuregs/_1376_ ),
    .A1(\soc/cpu/cpuregs/_1377_ ),
    .A2(\soc/cpu/cpuregs/_1378_ ),
    .A3(\soc/cpu/cpuregs/_1379_ ),
    .S0(\soc/cpu/cpuregs/_1025_ ),
    .S1(\soc/cpu/cpuregs/_1059_ ),
    .X(\soc/cpu/cpuregs/_1380_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2891_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1380_ ),
    .Y(\soc/cpu/cpuregs/_1381_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/cpuregs/_2892_  (.A(\soc/cpu/cpuregs/_1375_ ),
    .B(\soc/cpu/cpuregs/_1381_ ),
    .Y(\soc/cpu/cpuregs_rdata2[15] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2893_  (.A0(\soc/cpu/cpuregs/regs[16][16] ),
    .A1(\soc/cpu/cpuregs/regs[17][16] ),
    .A2(\soc/cpu/cpuregs/regs[20][16] ),
    .A3(\soc/cpu/cpuregs/regs[21][16] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1382_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2894_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1382_ ),
    .Y(\soc/cpu/cpuregs/_1383_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2895_  (.A0(\soc/cpu/cpuregs/regs[18][16] ),
    .A1(\soc/cpu/cpuregs/regs[19][16] ),
    .A2(\soc/cpu/cpuregs/regs[22][16] ),
    .A3(\soc/cpu/cpuregs/regs[23][16] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1384_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2896_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1384_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1385_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2897_  (.A0(\soc/cpu/cpuregs/regs[2][16] ),
    .A1(\soc/cpu/cpuregs/regs[3][16] ),
    .A2(\soc/cpu/cpuregs/regs[6][16] ),
    .A3(\soc/cpu/cpuregs/regs[7][16] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1386_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2898_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1386_ ),
    .Y(\soc/cpu/cpuregs/_1387_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2899_  (.A0(\soc/cpu/cpuregs/regs[0][16] ),
    .A1(\soc/cpu/cpuregs/regs[1][16] ),
    .A2(\soc/cpu/cpuregs/regs[4][16] ),
    .A3(\soc/cpu/cpuregs/regs[5][16] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1388_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2900_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1388_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1389_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2901_  (.A1(\soc/cpu/cpuregs/_1383_ ),
    .A2(\soc/cpu/cpuregs/_1385_ ),
    .B1(\soc/cpu/cpuregs/_1387_ ),
    .B2(\soc/cpu/cpuregs/_1389_ ),
    .Y(\soc/cpu/cpuregs/_1390_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2902_  (.A0(\soc/cpu/cpuregs/regs[24][16] ),
    .A1(\soc/cpu/cpuregs/regs[25][16] ),
    .A2(\soc/cpu/cpuregs/regs[28][16] ),
    .A3(\soc/cpu/cpuregs/regs[29][16] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1391_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2903_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1391_ ),
    .Y(\soc/cpu/cpuregs/_1392_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2904_  (.A0(\soc/cpu/cpuregs/regs[26][16] ),
    .A1(\soc/cpu/cpuregs/regs[27][16] ),
    .A2(\soc/cpu/cpuregs/regs[30][16] ),
    .A3(\soc/cpu/cpuregs/regs[31][16] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1393_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2905_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1393_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1394_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2906_  (.A0(\soc/cpu/cpuregs/regs[10][16] ),
    .A1(\soc/cpu/cpuregs/regs[11][16] ),
    .A2(\soc/cpu/cpuregs/regs[14][16] ),
    .A3(\soc/cpu/cpuregs/regs[15][16] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1395_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2907_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1395_ ),
    .Y(\soc/cpu/cpuregs/_1396_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2908_  (.A0(\soc/cpu/cpuregs/regs[8][16] ),
    .A1(\soc/cpu/cpuregs/regs[9][16] ),
    .A2(\soc/cpu/cpuregs/regs[12][16] ),
    .A3(\soc/cpu/cpuregs/regs[13][16] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1397_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2909_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1397_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1398_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_2910_  (.A1(\soc/cpu/cpuregs/_1392_ ),
    .A2(\soc/cpu/cpuregs/_1394_ ),
    .B1(\soc/cpu/cpuregs/_1396_ ),
    .B2(\soc/cpu/cpuregs/_1398_ ),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1399_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_2911_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1390_ ),
    .B1(\soc/cpu/cpuregs/_1399_ ),
    .X(\soc/cpu/cpuregs_rdata2[16] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2913_  (.A0(\soc/cpu/cpuregs/regs[2][17] ),
    .A1(\soc/cpu/cpuregs/regs[3][17] ),
    .A2(\soc/cpu/cpuregs/regs[6][17] ),
    .A3(\soc/cpu/cpuregs/regs[7][17] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1401_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2914_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1401_ ),
    .Y(\soc/cpu/cpuregs/_1402_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2915_  (.A0(\soc/cpu/cpuregs/regs[0][17] ),
    .A1(\soc/cpu/cpuregs/regs[1][17] ),
    .A2(\soc/cpu/cpuregs/regs[4][17] ),
    .A3(\soc/cpu/cpuregs/regs[5][17] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1403_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2916_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1403_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1404_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2917_  (.A0(\soc/cpu/cpuregs/regs[16][17] ),
    .A1(\soc/cpu/cpuregs/regs[17][17] ),
    .A2(\soc/cpu/cpuregs/regs[20][17] ),
    .A3(\soc/cpu/cpuregs/regs[21][17] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1405_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2918_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1405_ ),
    .Y(\soc/cpu/cpuregs/_1406_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2919_  (.A0(\soc/cpu/cpuregs/regs[18][17] ),
    .A1(\soc/cpu/cpuregs/regs[19][17] ),
    .A2(\soc/cpu/cpuregs/regs[22][17] ),
    .A3(\soc/cpu/cpuregs/regs[23][17] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1407_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2920_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1407_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1408_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2921_  (.A1(\soc/cpu/cpuregs/_1402_ ),
    .A2(\soc/cpu/cpuregs/_1404_ ),
    .B1(\soc/cpu/cpuregs/_1406_ ),
    .B2(\soc/cpu/cpuregs/_1408_ ),
    .Y(\soc/cpu/cpuregs/_1409_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2923_  (.A0(\soc/cpu/cpuregs/regs[10][17] ),
    .A1(\soc/cpu/cpuregs/regs[11][17] ),
    .A2(\soc/cpu/cpuregs/regs[14][17] ),
    .A3(\soc/cpu/cpuregs/regs[15][17] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1411_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2924_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1411_ ),
    .Y(\soc/cpu/cpuregs/_1412_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2925_  (.A0(\soc/cpu/cpuregs/regs[8][17] ),
    .A1(\soc/cpu/cpuregs/regs[9][17] ),
    .A2(\soc/cpu/cpuregs/regs[12][17] ),
    .A3(\soc/cpu/cpuregs/regs[13][17] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1413_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_2926_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1413_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1414_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2927_  (.A0(\soc/cpu/cpuregs/regs[24][17] ),
    .A1(\soc/cpu/cpuregs/regs[25][17] ),
    .A2(\soc/cpu/cpuregs/regs[28][17] ),
    .A3(\soc/cpu/cpuregs/regs[29][17] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1415_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2928_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1415_ ),
    .Y(\soc/cpu/cpuregs/_1416_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2929_  (.A0(\soc/cpu/cpuregs/regs[26][17] ),
    .A1(\soc/cpu/cpuregs/regs[27][17] ),
    .A2(\soc/cpu/cpuregs/regs[30][17] ),
    .A3(\soc/cpu/cpuregs/regs[31][17] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1417_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_2930_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1417_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1418_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_2932_  (.A1(\soc/cpu/cpuregs/_1412_ ),
    .A2(\soc/cpu/cpuregs/_1414_ ),
    .B1(\soc/cpu/cpuregs/_1416_ ),
    .B2(\soc/cpu/cpuregs/_1418_ ),
    .C1(net302),
    .Y(\soc/cpu/cpuregs/_1420_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2933_  (.A1(net302),
    .A2(\soc/cpu/cpuregs/_1409_ ),
    .B1(\soc/cpu/cpuregs/_1420_ ),
    .X(\soc/cpu/cpuregs_rdata2[17] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2934_  (.A0(\soc/cpu/cpuregs/regs[2][18] ),
    .A1(\soc/cpu/cpuregs/regs[3][18] ),
    .A2(\soc/cpu/cpuregs/regs[6][18] ),
    .A3(\soc/cpu/cpuregs/regs[7][18] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1421_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2935_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1421_ ),
    .Y(\soc/cpu/cpuregs/_1422_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2936_  (.A0(\soc/cpu/cpuregs/regs[0][18] ),
    .A1(\soc/cpu/cpuregs/regs[1][18] ),
    .A2(\soc/cpu/cpuregs/regs[4][18] ),
    .A3(\soc/cpu/cpuregs/regs[5][18] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1423_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2937_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1423_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1424_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2938_  (.A0(\soc/cpu/cpuregs/regs[18][18] ),
    .A1(\soc/cpu/cpuregs/regs[19][18] ),
    .A2(\soc/cpu/cpuregs/regs[22][18] ),
    .A3(\soc/cpu/cpuregs/regs[23][18] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1425_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2939_  (.A0(\soc/cpu/cpuregs/regs[16][18] ),
    .A1(\soc/cpu/cpuregs/regs[17][18] ),
    .A2(\soc/cpu/cpuregs/regs[20][18] ),
    .A3(\soc/cpu/cpuregs/regs[21][18] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1426_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2940_  (.A0(\soc/cpu/cpuregs/_1425_ ),
    .A1(\soc/cpu/cpuregs/_1426_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1427_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_2941_  (.A1(\soc/cpu/cpuregs/_1422_ ),
    .A2(\soc/cpu/cpuregs/_1424_ ),
    .B1(\soc/cpu/cpuregs/_1427_ ),
    .B2(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1428_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2942_  (.A0(\soc/cpu/cpuregs/regs[26][18] ),
    .A1(\soc/cpu/cpuregs/regs[27][18] ),
    .A2(\soc/cpu/cpuregs/regs[30][18] ),
    .A3(\soc/cpu/cpuregs/regs[31][18] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1429_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2943_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1429_ ),
    .Y(\soc/cpu/cpuregs/_1430_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2944_  (.A0(\soc/cpu/cpuregs/regs[24][18] ),
    .A1(\soc/cpu/cpuregs/regs[25][18] ),
    .A2(\soc/cpu/cpuregs/regs[28][18] ),
    .A3(\soc/cpu/cpuregs/regs[29][18] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1431_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2945_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1431_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1432_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2946_  (.A0(\soc/cpu/cpuregs/regs[10][18] ),
    .A1(\soc/cpu/cpuregs/regs[11][18] ),
    .A2(\soc/cpu/cpuregs/regs[14][18] ),
    .A3(\soc/cpu/cpuregs/regs[15][18] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1433_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2947_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1433_ ),
    .Y(\soc/cpu/cpuregs/_1434_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2948_  (.A0(\soc/cpu/cpuregs/regs[8][18] ),
    .A1(\soc/cpu/cpuregs/regs[9][18] ),
    .A2(\soc/cpu/cpuregs/regs[12][18] ),
    .A3(\soc/cpu/cpuregs/regs[13][18] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1435_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2949_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1435_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1436_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2950_  (.A1(\soc/cpu/cpuregs/_1430_ ),
    .A2(\soc/cpu/cpuregs/_1432_ ),
    .B1(\soc/cpu/cpuregs/_1434_ ),
    .B2(\soc/cpu/cpuregs/_1436_ ),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1437_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2951_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1428_ ),
    .B1(\soc/cpu/cpuregs/_1437_ ),
    .X(\soc/cpu/cpuregs_rdata2[18] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2953_  (.A0(\soc/cpu/cpuregs/regs[2][19] ),
    .A1(\soc/cpu/cpuregs/regs[3][19] ),
    .A2(\soc/cpu/cpuregs/regs[6][19] ),
    .A3(\soc/cpu/cpuregs/regs[7][19] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1439_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2954_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1439_ ),
    .Y(\soc/cpu/cpuregs/_1440_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2955_  (.A0(\soc/cpu/cpuregs/regs[0][19] ),
    .A1(\soc/cpu/cpuregs/regs[1][19] ),
    .A2(\soc/cpu/cpuregs/regs[4][19] ),
    .A3(\soc/cpu/cpuregs/regs[5][19] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1441_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_2956_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1441_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1442_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2958_  (.A0(\soc/cpu/cpuregs/regs[16][19] ),
    .A1(\soc/cpu/cpuregs/regs[17][19] ),
    .A2(\soc/cpu/cpuregs/regs[20][19] ),
    .A3(\soc/cpu/cpuregs/regs[21][19] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1444_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2959_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1444_ ),
    .Y(\soc/cpu/cpuregs/_1445_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2960_  (.A0(\soc/cpu/cpuregs/regs[18][19] ),
    .A1(\soc/cpu/cpuregs/regs[19][19] ),
    .A2(\soc/cpu/cpuregs/regs[22][19] ),
    .A3(\soc/cpu/cpuregs/regs[23][19] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1446_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_2961_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1446_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1447_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/cpuregs/_2962_  (.A1(\soc/cpu/cpuregs/_1440_ ),
    .A2(\soc/cpu/cpuregs/_1442_ ),
    .B1(\soc/cpu/cpuregs/_1445_ ),
    .B2(\soc/cpu/cpuregs/_1447_ ),
    .Y(\soc/cpu/cpuregs/_1448_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2964_  (.A0(\soc/cpu/cpuregs/regs[10][19] ),
    .A1(\soc/cpu/cpuregs/regs[11][19] ),
    .A2(\soc/cpu/cpuregs/regs[14][19] ),
    .A3(\soc/cpu/cpuregs/regs[15][19] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1450_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2965_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1450_ ),
    .Y(\soc/cpu/cpuregs/_1451_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2966_  (.A0(\soc/cpu/cpuregs/regs[8][19] ),
    .A1(\soc/cpu/cpuregs/regs[9][19] ),
    .A2(\soc/cpu/cpuregs/regs[12][19] ),
    .A3(\soc/cpu/cpuregs/regs[13][19] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1452_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2967_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1452_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1453_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2968_  (.A0(\soc/cpu/cpuregs/regs[24][19] ),
    .A1(\soc/cpu/cpuregs/regs[25][19] ),
    .A2(\soc/cpu/cpuregs/regs[28][19] ),
    .A3(\soc/cpu/cpuregs/regs[29][19] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1454_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2969_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1454_ ),
    .Y(\soc/cpu/cpuregs/_1455_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2970_  (.A0(\soc/cpu/cpuregs/regs[26][19] ),
    .A1(\soc/cpu/cpuregs/regs[27][19] ),
    .A2(\soc/cpu/cpuregs/regs[30][19] ),
    .A3(\soc/cpu/cpuregs/regs[31][19] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1456_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2971_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1456_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1457_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2972_  (.A1(\soc/cpu/cpuregs/_1451_ ),
    .A2(\soc/cpu/cpuregs/_1453_ ),
    .B1(\soc/cpu/cpuregs/_1455_ ),
    .B2(\soc/cpu/cpuregs/_1457_ ),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1458_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2973_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1448_ ),
    .B1(\soc/cpu/cpuregs/_1458_ ),
    .X(\soc/cpu/cpuregs_rdata2[19] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2974_  (.A0(\soc/cpu/cpuregs/regs[16][20] ),
    .A1(\soc/cpu/cpuregs/regs[17][20] ),
    .A2(\soc/cpu/cpuregs/regs[20][20] ),
    .A3(\soc/cpu/cpuregs/regs[21][20] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1459_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2975_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1459_ ),
    .Y(\soc/cpu/cpuregs/_1460_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2976_  (.A0(\soc/cpu/cpuregs/regs[18][20] ),
    .A1(\soc/cpu/cpuregs/regs[19][20] ),
    .A2(\soc/cpu/cpuregs/regs[22][20] ),
    .A3(\soc/cpu/cpuregs/regs[23][20] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1461_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2977_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1461_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1462_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2978_  (.A0(\soc/cpu/cpuregs/regs[2][20] ),
    .A1(\soc/cpu/cpuregs/regs[3][20] ),
    .A2(\soc/cpu/cpuregs/regs[6][20] ),
    .A3(\soc/cpu/cpuregs/regs[7][20] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1463_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2979_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1463_ ),
    .Y(\soc/cpu/cpuregs/_1464_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2980_  (.A0(\soc/cpu/cpuregs/regs[0][20] ),
    .A1(\soc/cpu/cpuregs/regs[1][20] ),
    .A2(\soc/cpu/cpuregs/regs[4][20] ),
    .A3(\soc/cpu/cpuregs/regs[5][20] ),
    .S0(net318),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1465_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_2981_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1465_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1466_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_2982_  (.A1(\soc/cpu/cpuregs/_1460_ ),
    .A2(\soc/cpu/cpuregs/_1462_ ),
    .B1(\soc/cpu/cpuregs/_1464_ ),
    .B2(\soc/cpu/cpuregs/_1466_ ),
    .Y(\soc/cpu/cpuregs/_1467_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2983_  (.A0(\soc/cpu/cpuregs/regs[24][20] ),
    .A1(\soc/cpu/cpuregs/regs[25][20] ),
    .A2(\soc/cpu/cpuregs/regs[28][20] ),
    .A3(\soc/cpu/cpuregs/regs[29][20] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1468_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_2984_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1468_ ),
    .Y(\soc/cpu/cpuregs/_1469_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2985_  (.A0(\soc/cpu/cpuregs/regs[26][20] ),
    .A1(\soc/cpu/cpuregs/regs[27][20] ),
    .A2(\soc/cpu/cpuregs/regs[30][20] ),
    .A3(\soc/cpu/cpuregs/regs[31][20] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1470_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_2986_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1470_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1471_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2987_  (.A0(\soc/cpu/cpuregs/regs[10][20] ),
    .A1(\soc/cpu/cpuregs/regs[11][20] ),
    .A2(\soc/cpu/cpuregs/regs[14][20] ),
    .A3(\soc/cpu/cpuregs/regs[15][20] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1472_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2988_  (.A0(\soc/cpu/cpuregs/regs[8][20] ),
    .A1(\soc/cpu/cpuregs/regs[9][20] ),
    .A2(\soc/cpu/cpuregs/regs[12][20] ),
    .A3(\soc/cpu/cpuregs/regs[13][20] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1473_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_2989_  (.A0(\soc/cpu/cpuregs/_1472_ ),
    .A1(\soc/cpu/cpuregs/_1473_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1474_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_2990_  (.A1(\soc/cpu/cpuregs/_1469_ ),
    .A2(\soc/cpu/cpuregs/_1471_ ),
    .B1(\soc/cpu/cpuregs/_1474_ ),
    .B2(net299),
    .C1(net302),
    .Y(\soc/cpu/cpuregs/_1475_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_2991_  (.A1(net302),
    .A2(\soc/cpu/cpuregs/_1467_ ),
    .B1(\soc/cpu/cpuregs/_1475_ ),
    .X(\soc/cpu/cpuregs_rdata2[20] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2992_  (.A0(\soc/cpu/cpuregs/regs[2][21] ),
    .A1(\soc/cpu/cpuregs/regs[3][21] ),
    .A2(\soc/cpu/cpuregs/regs[6][21] ),
    .A3(\soc/cpu/cpuregs/regs[7][21] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1476_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2993_  (.A0(\soc/cpu/cpuregs/regs[0][21] ),
    .A1(\soc/cpu/cpuregs/regs[1][21] ),
    .A2(\soc/cpu/cpuregs/regs[4][21] ),
    .A3(\soc/cpu/cpuregs/regs[5][21] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1477_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_2994_  (.A0(\soc/cpu/cpuregs/_1476_ ),
    .A1(\soc/cpu/cpuregs/_1477_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1478_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2995_  (.A0(\soc/cpu/cpuregs/regs[18][21] ),
    .A1(\soc/cpu/cpuregs/regs[19][21] ),
    .A2(\soc/cpu/cpuregs/regs[22][21] ),
    .A3(\soc/cpu/cpuregs/regs[23][21] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1479_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_2996_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1479_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1480_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_2997_  (.A0(\soc/cpu/cpuregs/regs[16][21] ),
    .A1(\soc/cpu/cpuregs/regs[17][21] ),
    .A2(\soc/cpu/cpuregs/regs[20][21] ),
    .A3(\soc/cpu/cpuregs/regs[21][21] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1481_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_2998_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1481_ ),
    .Y(\soc/cpu/cpuregs/_1482_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/cpu/cpuregs/_2999_  (.A1(\soc/cpu/cpuregs/_1059_ ),
    .A2(\soc/cpu/cpuregs/_1478_ ),
    .B1(\soc/cpu/cpuregs/_1480_ ),
    .B2(\soc/cpu/cpuregs/_1482_ ),
    .Y(\soc/cpu/cpuregs/_1483_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3000_  (.A0(\soc/cpu/cpuregs/regs[10][21] ),
    .A1(\soc/cpu/cpuregs/regs[11][21] ),
    .A2(\soc/cpu/cpuregs/regs[14][21] ),
    .A3(\soc/cpu/cpuregs/regs[15][21] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1484_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3001_  (.A0(\soc/cpu/cpuregs/regs[8][21] ),
    .A1(\soc/cpu/cpuregs/regs[9][21] ),
    .A2(\soc/cpu/cpuregs/regs[12][21] ),
    .A3(\soc/cpu/cpuregs/regs[13][21] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1485_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3002_  (.A0(\soc/cpu/cpuregs/_1484_ ),
    .A1(\soc/cpu/cpuregs/_1485_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1486_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3003_  (.A0(\soc/cpu/cpuregs/regs[26][21] ),
    .A1(\soc/cpu/cpuregs/regs[27][21] ),
    .A2(\soc/cpu/cpuregs/regs[30][21] ),
    .A3(\soc/cpu/cpuregs/regs[31][21] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1487_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3004_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1487_ ),
    .Y(\soc/cpu/cpuregs/_1488_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3005_  (.A0(\soc/cpu/cpuregs/regs[24][21] ),
    .A1(\soc/cpu/cpuregs/regs[25][21] ),
    .A2(\soc/cpu/cpuregs/regs[28][21] ),
    .A3(\soc/cpu/cpuregs/regs[29][21] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1489_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3006_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1489_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1490_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3007_  (.A1(net300),
    .A2(\soc/cpu/cpuregs/_1486_ ),
    .B1(\soc/cpu/cpuregs/_1488_ ),
    .B2(\soc/cpu/cpuregs/_1490_ ),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1491_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3008_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1483_ ),
    .B1(\soc/cpu/cpuregs/_1491_ ),
    .X(\soc/cpu/cpuregs_rdata2[21] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3009_  (.A0(\soc/cpu/cpuregs/regs[2][22] ),
    .A1(\soc/cpu/cpuregs/regs[3][22] ),
    .A2(\soc/cpu/cpuregs/regs[6][22] ),
    .A3(\soc/cpu/cpuregs/regs[7][22] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1492_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3010_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1492_ ),
    .Y(\soc/cpu/cpuregs/_1493_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3011_  (.A0(\soc/cpu/cpuregs/regs[0][22] ),
    .A1(\soc/cpu/cpuregs/regs[1][22] ),
    .A2(\soc/cpu/cpuregs/regs[4][22] ),
    .A3(\soc/cpu/cpuregs/regs[5][22] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1494_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3012_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1494_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1495_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3013_  (.A0(\soc/cpu/cpuregs/regs[16][22] ),
    .A1(\soc/cpu/cpuregs/regs[17][22] ),
    .A2(\soc/cpu/cpuregs/regs[20][22] ),
    .A3(\soc/cpu/cpuregs/regs[21][22] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1496_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3014_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1496_ ),
    .Y(\soc/cpu/cpuregs/_1497_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3015_  (.A0(\soc/cpu/cpuregs/regs[18][22] ),
    .A1(\soc/cpu/cpuregs/regs[19][22] ),
    .A2(\soc/cpu/cpuregs/regs[22][22] ),
    .A3(\soc/cpu/cpuregs/regs[23][22] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1498_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3016_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1498_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1499_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3017_  (.A1(\soc/cpu/cpuregs/_1493_ ),
    .A2(\soc/cpu/cpuregs/_1495_ ),
    .B1(\soc/cpu/cpuregs/_1497_ ),
    .B2(\soc/cpu/cpuregs/_1499_ ),
    .Y(\soc/cpu/cpuregs/_1500_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3018_  (.A0(\soc/cpu/cpuregs/regs[10][22] ),
    .A1(\soc/cpu/cpuregs/regs[11][22] ),
    .A2(\soc/cpu/cpuregs/regs[14][22] ),
    .A3(\soc/cpu/cpuregs/regs[15][22] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1501_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3019_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1501_ ),
    .Y(\soc/cpu/cpuregs/_1502_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3020_  (.A0(\soc/cpu/cpuregs/regs[8][22] ),
    .A1(\soc/cpu/cpuregs/regs[9][22] ),
    .A2(\soc/cpu/cpuregs/regs[12][22] ),
    .A3(\soc/cpu/cpuregs/regs[13][22] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1503_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3021_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1503_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1504_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3022_  (.A0(\soc/cpu/cpuregs/regs[24][22] ),
    .A1(\soc/cpu/cpuregs/regs[25][22] ),
    .A2(\soc/cpu/cpuregs/regs[28][22] ),
    .A3(\soc/cpu/cpuregs/regs[29][22] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1505_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3023_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1505_ ),
    .Y(\soc/cpu/cpuregs/_1506_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3024_  (.A0(\soc/cpu/cpuregs/regs[26][22] ),
    .A1(\soc/cpu/cpuregs/regs[27][22] ),
    .A2(\soc/cpu/cpuregs/regs[30][22] ),
    .A3(\soc/cpu/cpuregs/regs[31][22] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1507_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3025_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1507_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1508_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3026_  (.A1(\soc/cpu/cpuregs/_1502_ ),
    .A2(\soc/cpu/cpuregs/_1504_ ),
    .B1(\soc/cpu/cpuregs/_1506_ ),
    .B2(\soc/cpu/cpuregs/_1508_ ),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1509_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3027_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1500_ ),
    .B1(\soc/cpu/cpuregs/_1509_ ),
    .X(\soc/cpu/cpuregs_rdata2[22] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3028_  (.A0(\soc/cpu/cpuregs/regs[16][23] ),
    .A1(\soc/cpu/cpuregs/regs[17][23] ),
    .A2(\soc/cpu/cpuregs/regs[20][23] ),
    .A3(\soc/cpu/cpuregs/regs[21][23] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1510_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3029_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1510_ ),
    .Y(\soc/cpu/cpuregs/_1511_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3030_  (.A0(\soc/cpu/cpuregs/regs[18][23] ),
    .A1(\soc/cpu/cpuregs/regs[19][23] ),
    .A2(\soc/cpu/cpuregs/regs[22][23] ),
    .A3(\soc/cpu/cpuregs/regs[23][23] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1512_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3031_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1512_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1513_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3032_  (.A0(\soc/cpu/cpuregs/regs[2][23] ),
    .A1(\soc/cpu/cpuregs/regs[3][23] ),
    .A2(\soc/cpu/cpuregs/regs[6][23] ),
    .A3(\soc/cpu/cpuregs/regs[7][23] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1514_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3033_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1514_ ),
    .Y(\soc/cpu/cpuregs/_1515_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3034_  (.A0(\soc/cpu/cpuregs/regs[0][23] ),
    .A1(\soc/cpu/cpuregs/regs[1][23] ),
    .A2(\soc/cpu/cpuregs/regs[4][23] ),
    .A3(\soc/cpu/cpuregs/regs[5][23] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1516_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3035_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1516_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1517_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3036_  (.A1(\soc/cpu/cpuregs/_1511_ ),
    .A2(\soc/cpu/cpuregs/_1513_ ),
    .B1(\soc/cpu/cpuregs/_1515_ ),
    .B2(\soc/cpu/cpuregs/_1517_ ),
    .Y(\soc/cpu/cpuregs/_1518_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3037_  (.A0(\soc/cpu/cpuregs/regs[24][23] ),
    .A1(\soc/cpu/cpuregs/regs[25][23] ),
    .A2(\soc/cpu/cpuregs/regs[28][23] ),
    .A3(\soc/cpu/cpuregs/regs[29][23] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1519_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3038_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1519_ ),
    .Y(\soc/cpu/cpuregs/_1520_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3039_  (.A0(\soc/cpu/cpuregs/regs[26][23] ),
    .A1(\soc/cpu/cpuregs/regs[27][23] ),
    .A2(\soc/cpu/cpuregs/regs[30][23] ),
    .A3(\soc/cpu/cpuregs/regs[31][23] ),
    .S0(net317),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1521_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3040_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1521_ ),
    .B1(net298),
    .Y(\soc/cpu/cpuregs/_1522_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3041_  (.A0(\soc/cpu/cpuregs/regs[10][23] ),
    .A1(\soc/cpu/cpuregs/regs[11][23] ),
    .A2(\soc/cpu/cpuregs/regs[14][23] ),
    .A3(\soc/cpu/cpuregs/regs[15][23] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1523_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3042_  (.A0(\soc/cpu/cpuregs/regs[8][23] ),
    .A1(\soc/cpu/cpuregs/regs[9][23] ),
    .A2(\soc/cpu/cpuregs/regs[12][23] ),
    .A3(\soc/cpu/cpuregs/regs[13][23] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1524_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_3043_  (.A0(\soc/cpu/cpuregs/_1523_ ),
    .A1(\soc/cpu/cpuregs/_1524_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1525_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3044_  (.A1(\soc/cpu/cpuregs/_1520_ ),
    .A2(\soc/cpu/cpuregs/_1522_ ),
    .B1(\soc/cpu/cpuregs/_1525_ ),
    .B2(net298),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1526_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3045_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1518_ ),
    .B1(\soc/cpu/cpuregs/_1526_ ),
    .X(\soc/cpu/cpuregs_rdata2[23] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3046_  (.A0(\soc/cpu/cpuregs/regs[16][24] ),
    .A1(\soc/cpu/cpuregs/regs[17][24] ),
    .A2(\soc/cpu/cpuregs/regs[20][24] ),
    .A3(\soc/cpu/cpuregs/regs[21][24] ),
    .S0(net326),
    .S1(\soc/cpu/cpuregs_raddr2[2] ),
    .X(\soc/cpu/cpuregs/_1527_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3047_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1527_ ),
    .Y(\soc/cpu/cpuregs/_1528_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3048_  (.A0(\soc/cpu/cpuregs/regs[18][24] ),
    .A1(\soc/cpu/cpuregs/regs[19][24] ),
    .A2(\soc/cpu/cpuregs/regs[22][24] ),
    .A3(\soc/cpu/cpuregs/regs[23][24] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1529_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3049_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1529_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1530_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3050_  (.A0(\soc/cpu/cpuregs/regs[2][24] ),
    .A1(\soc/cpu/cpuregs/regs[3][24] ),
    .A2(\soc/cpu/cpuregs/regs[6][24] ),
    .A3(\soc/cpu/cpuregs/regs[7][24] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1531_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3051_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1531_ ),
    .Y(\soc/cpu/cpuregs/_1532_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3052_  (.A0(\soc/cpu/cpuregs/regs[0][24] ),
    .A1(\soc/cpu/cpuregs/regs[1][24] ),
    .A2(\soc/cpu/cpuregs/regs[4][24] ),
    .A3(\soc/cpu/cpuregs/regs[5][24] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1533_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3053_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1533_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1534_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3054_  (.A1(\soc/cpu/cpuregs/_1528_ ),
    .A2(\soc/cpu/cpuregs/_1530_ ),
    .B1(\soc/cpu/cpuregs/_1532_ ),
    .B2(\soc/cpu/cpuregs/_1534_ ),
    .Y(\soc/cpu/cpuregs/_1535_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3055_  (.A0(\soc/cpu/cpuregs/regs[24][24] ),
    .A1(\soc/cpu/cpuregs/regs[25][24] ),
    .A2(\soc/cpu/cpuregs/regs[28][24] ),
    .A3(\soc/cpu/cpuregs/regs[29][24] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1536_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3056_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1536_ ),
    .Y(\soc/cpu/cpuregs/_1537_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3057_  (.A0(\soc/cpu/cpuregs/regs[26][24] ),
    .A1(\soc/cpu/cpuregs/regs[27][24] ),
    .A2(\soc/cpu/cpuregs/regs[30][24] ),
    .A3(\soc/cpu/cpuregs/regs[31][24] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1538_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3058_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1538_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1539_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3059_  (.A0(\soc/cpu/cpuregs/regs[10][24] ),
    .A1(\soc/cpu/cpuregs/regs[11][24] ),
    .A2(\soc/cpu/cpuregs/regs[14][24] ),
    .A3(\soc/cpu/cpuregs/regs[15][24] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1540_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3060_  (.A0(\soc/cpu/cpuregs/regs[8][24] ),
    .A1(\soc/cpu/cpuregs/regs[9][24] ),
    .A2(\soc/cpu/cpuregs/regs[12][24] ),
    .A3(\soc/cpu/cpuregs/regs[13][24] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1541_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3061_  (.A0(\soc/cpu/cpuregs/_1540_ ),
    .A1(\soc/cpu/cpuregs/_1541_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1542_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3062_  (.A1(\soc/cpu/cpuregs/_1537_ ),
    .A2(\soc/cpu/cpuregs/_1539_ ),
    .B1(\soc/cpu/cpuregs/_1542_ ),
    .B2(net301),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1543_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3063_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1535_ ),
    .B1(\soc/cpu/cpuregs/_1543_ ),
    .X(\soc/cpu/cpuregs_rdata2[24] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3064_  (.A0(\soc/cpu/cpuregs/regs[16][25] ),
    .A1(\soc/cpu/cpuregs/regs[17][25] ),
    .A2(\soc/cpu/cpuregs/regs[20][25] ),
    .A3(\soc/cpu/cpuregs/regs[21][25] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1544_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3065_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1544_ ),
    .Y(\soc/cpu/cpuregs/_1545_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3066_  (.A0(\soc/cpu/cpuregs/regs[18][25] ),
    .A1(\soc/cpu/cpuregs/regs[19][25] ),
    .A2(\soc/cpu/cpuregs/regs[22][25] ),
    .A3(\soc/cpu/cpuregs/regs[23][25] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1546_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3067_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1546_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1547_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3068_  (.A0(\soc/cpu/cpuregs/regs[2][25] ),
    .A1(\soc/cpu/cpuregs/regs[3][25] ),
    .A2(\soc/cpu/cpuregs/regs[6][25] ),
    .A3(\soc/cpu/cpuregs/regs[7][25] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1548_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3069_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1548_ ),
    .Y(\soc/cpu/cpuregs/_1549_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3070_  (.A0(\soc/cpu/cpuregs/regs[0][25] ),
    .A1(\soc/cpu/cpuregs/regs[1][25] ),
    .A2(\soc/cpu/cpuregs/regs[4][25] ),
    .A3(\soc/cpu/cpuregs/regs[5][25] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1550_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3071_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1550_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1551_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3072_  (.A1(\soc/cpu/cpuregs/_1545_ ),
    .A2(\soc/cpu/cpuregs/_1547_ ),
    .B1(\soc/cpu/cpuregs/_1549_ ),
    .B2(\soc/cpu/cpuregs/_1551_ ),
    .Y(\soc/cpu/cpuregs/_1552_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3073_  (.A0(\soc/cpu/cpuregs/regs[24][25] ),
    .A1(\soc/cpu/cpuregs/regs[25][25] ),
    .A2(\soc/cpu/cpuregs/regs[28][25] ),
    .A3(\soc/cpu/cpuregs/regs[29][25] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1553_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3074_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1553_ ),
    .Y(\soc/cpu/cpuregs/_1554_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3075_  (.A0(\soc/cpu/cpuregs/regs[26][25] ),
    .A1(\soc/cpu/cpuregs/regs[27][25] ),
    .A2(\soc/cpu/cpuregs/regs[30][25] ),
    .A3(\soc/cpu/cpuregs/regs[31][25] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1555_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3076_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1555_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1556_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3077_  (.A0(\soc/cpu/cpuregs/regs[10][25] ),
    .A1(\soc/cpu/cpuregs/regs[11][25] ),
    .A2(\soc/cpu/cpuregs/regs[14][25] ),
    .A3(\soc/cpu/cpuregs/regs[15][25] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1557_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3078_  (.A0(\soc/cpu/cpuregs/regs[8][25] ),
    .A1(\soc/cpu/cpuregs/regs[9][25] ),
    .A2(\soc/cpu/cpuregs/regs[12][25] ),
    .A3(\soc/cpu/cpuregs/regs[13][25] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1558_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3079_  (.A0(\soc/cpu/cpuregs/_1557_ ),
    .A1(\soc/cpu/cpuregs/_1558_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1559_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3080_  (.A1(\soc/cpu/cpuregs/_1554_ ),
    .A2(\soc/cpu/cpuregs/_1556_ ),
    .B1(\soc/cpu/cpuregs/_1559_ ),
    .B2(net299),
    .C1(net302),
    .Y(\soc/cpu/cpuregs/_1560_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3081_  (.A1(net302),
    .A2(\soc/cpu/cpuregs/_1552_ ),
    .B1(\soc/cpu/cpuregs/_1560_ ),
    .X(\soc/cpu/cpuregs_rdata2[25] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3082_  (.A0(\soc/cpu/cpuregs/regs[2][26] ),
    .A1(\soc/cpu/cpuregs/regs[3][26] ),
    .A2(\soc/cpu/cpuregs/regs[6][26] ),
    .A3(\soc/cpu/cpuregs/regs[7][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1561_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3083_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1561_ ),
    .Y(\soc/cpu/cpuregs/_1562_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3084_  (.A0(\soc/cpu/cpuregs/regs[0][26] ),
    .A1(\soc/cpu/cpuregs/regs[1][26] ),
    .A2(\soc/cpu/cpuregs/regs[4][26] ),
    .A3(\soc/cpu/cpuregs/regs[5][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1563_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3085_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1563_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1564_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3086_  (.A0(\soc/cpu/cpuregs/regs[16][26] ),
    .A1(\soc/cpu/cpuregs/regs[17][26] ),
    .A2(\soc/cpu/cpuregs/regs[20][26] ),
    .A3(\soc/cpu/cpuregs/regs[21][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1565_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3087_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1565_ ),
    .Y(\soc/cpu/cpuregs/_1566_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3088_  (.A0(\soc/cpu/cpuregs/regs[18][26] ),
    .A1(\soc/cpu/cpuregs/regs[19][26] ),
    .A2(\soc/cpu/cpuregs/regs[22][26] ),
    .A3(\soc/cpu/cpuregs/regs[23][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1567_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3089_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1567_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1568_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3090_  (.A1(\soc/cpu/cpuregs/_1562_ ),
    .A2(\soc/cpu/cpuregs/_1564_ ),
    .B1(\soc/cpu/cpuregs/_1566_ ),
    .B2(\soc/cpu/cpuregs/_1568_ ),
    .Y(\soc/cpu/cpuregs/_1569_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3091_  (.A0(\soc/cpu/cpuregs/regs[10][26] ),
    .A1(\soc/cpu/cpuregs/regs[11][26] ),
    .A2(\soc/cpu/cpuregs/regs[14][26] ),
    .A3(\soc/cpu/cpuregs/regs[15][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1570_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3092_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1570_ ),
    .Y(\soc/cpu/cpuregs/_1571_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3093_  (.A0(\soc/cpu/cpuregs/regs[8][26] ),
    .A1(\soc/cpu/cpuregs/regs[9][26] ),
    .A2(\soc/cpu/cpuregs/regs[12][26] ),
    .A3(\soc/cpu/cpuregs/regs[13][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1572_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3094_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1572_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1573_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3095_  (.A0(\soc/cpu/cpuregs/regs[24][26] ),
    .A1(\soc/cpu/cpuregs/regs[25][26] ),
    .A2(\soc/cpu/cpuregs/regs[28][26] ),
    .A3(\soc/cpu/cpuregs/regs[29][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1574_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3096_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1574_ ),
    .Y(\soc/cpu/cpuregs/_1575_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3097_  (.A0(\soc/cpu/cpuregs/regs[26][26] ),
    .A1(\soc/cpu/cpuregs/regs[27][26] ),
    .A2(\soc/cpu/cpuregs/regs[30][26] ),
    .A3(\soc/cpu/cpuregs/regs[31][26] ),
    .S0(net321),
    .S1(net308),
    .X(\soc/cpu/cpuregs/_1576_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3098_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1576_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1577_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3099_  (.A1(\soc/cpu/cpuregs/_1571_ ),
    .A2(\soc/cpu/cpuregs/_1573_ ),
    .B1(\soc/cpu/cpuregs/_1575_ ),
    .B2(\soc/cpu/cpuregs/_1577_ ),
    .C1(net304),
    .Y(\soc/cpu/cpuregs/_1578_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/cpuregs/_3100_  (.A1(net304),
    .A2(\soc/cpu/cpuregs/_1569_ ),
    .B1(\soc/cpu/cpuregs/_1578_ ),
    .X(\soc/cpu/cpuregs_rdata2[26] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3101_  (.A0(\soc/cpu/cpuregs/regs[16][27] ),
    .A1(\soc/cpu/cpuregs/regs[17][27] ),
    .A2(\soc/cpu/cpuregs/regs[20][27] ),
    .A3(\soc/cpu/cpuregs/regs[21][27] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1579_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3102_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1579_ ),
    .Y(\soc/cpu/cpuregs/_1580_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3103_  (.A0(\soc/cpu/cpuregs/regs[18][27] ),
    .A1(\soc/cpu/cpuregs/regs[19][27] ),
    .A2(\soc/cpu/cpuregs/regs[22][27] ),
    .A3(\soc/cpu/cpuregs/regs[23][27] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1581_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3104_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1581_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1582_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3105_  (.A0(\soc/cpu/cpuregs/regs[2][27] ),
    .A1(\soc/cpu/cpuregs/regs[3][27] ),
    .A2(\soc/cpu/cpuregs/regs[6][27] ),
    .A3(\soc/cpu/cpuregs/regs[7][27] ),
    .S0(net320),
    .S1(net306),
    .X(\soc/cpu/cpuregs/_1583_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3106_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1583_ ),
    .Y(\soc/cpu/cpuregs/_1584_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3107_  (.A0(\soc/cpu/cpuregs/regs[0][27] ),
    .A1(\soc/cpu/cpuregs/regs[1][27] ),
    .A2(\soc/cpu/cpuregs/regs[4][27] ),
    .A3(\soc/cpu/cpuregs/regs[5][27] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1585_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3108_  (.A1(net313),
    .A2(\soc/cpu/cpuregs/_1585_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1586_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3109_  (.A1(\soc/cpu/cpuregs/_1580_ ),
    .A2(\soc/cpu/cpuregs/_1582_ ),
    .B1(\soc/cpu/cpuregs/_1584_ ),
    .B2(\soc/cpu/cpuregs/_1586_ ),
    .Y(\soc/cpu/cpuregs/_1587_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3110_  (.A0(\soc/cpu/cpuregs/regs[24][27] ),
    .A1(\soc/cpu/cpuregs/regs[25][27] ),
    .A2(\soc/cpu/cpuregs/regs[28][27] ),
    .A3(\soc/cpu/cpuregs/regs[29][27] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1588_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3111_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1588_ ),
    .Y(\soc/cpu/cpuregs/_1589_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3112_  (.A0(\soc/cpu/cpuregs/regs[26][27] ),
    .A1(\soc/cpu/cpuregs/regs[27][27] ),
    .A2(\soc/cpu/cpuregs/regs[30][27] ),
    .A3(\soc/cpu/cpuregs/regs[31][27] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1590_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3113_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1590_ ),
    .B1(net299),
    .Y(\soc/cpu/cpuregs/_1591_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3114_  (.A0(\soc/cpu/cpuregs/regs[10][27] ),
    .A1(\soc/cpu/cpuregs/regs[11][27] ),
    .A2(\soc/cpu/cpuregs/regs[14][27] ),
    .A3(\soc/cpu/cpuregs/regs[15][27] ),
    .S0(net316),
    .S1(net305),
    .X(\soc/cpu/cpuregs/_1592_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3115_  (.A0(\soc/cpu/cpuregs/regs[8][27] ),
    .A1(\soc/cpu/cpuregs/regs[9][27] ),
    .A2(\soc/cpu/cpuregs/regs[12][27] ),
    .A3(\soc/cpu/cpuregs/regs[13][27] ),
    .S0(net319),
    .S1(net307),
    .X(\soc/cpu/cpuregs/_1593_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3116_  (.A0(\soc/cpu/cpuregs/_1592_ ),
    .A1(\soc/cpu/cpuregs/_1593_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1594_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3117_  (.A1(\soc/cpu/cpuregs/_1589_ ),
    .A2(\soc/cpu/cpuregs/_1591_ ),
    .B1(\soc/cpu/cpuregs/_1594_ ),
    .B2(net299),
    .C1(net302),
    .Y(\soc/cpu/cpuregs/_1595_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3118_  (.A1(net302),
    .A2(\soc/cpu/cpuregs/_1587_ ),
    .B1(\soc/cpu/cpuregs/_1595_ ),
    .X(\soc/cpu/cpuregs_rdata2[27] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3119_  (.A0(\soc/cpu/cpuregs/regs[16][28] ),
    .A1(\soc/cpu/cpuregs/regs[17][28] ),
    .A2(\soc/cpu/cpuregs/regs[20][28] ),
    .A3(\soc/cpu/cpuregs/regs[21][28] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1596_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3120_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1596_ ),
    .Y(\soc/cpu/cpuregs/_1597_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3121_  (.A0(\soc/cpu/cpuregs/regs[18][28] ),
    .A1(\soc/cpu/cpuregs/regs[19][28] ),
    .A2(\soc/cpu/cpuregs/regs[22][28] ),
    .A3(\soc/cpu/cpuregs/regs[23][28] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1598_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3122_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1598_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1599_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3123_  (.A0(\soc/cpu/cpuregs/regs[2][28] ),
    .A1(\soc/cpu/cpuregs/regs[3][28] ),
    .A2(\soc/cpu/cpuregs/regs[6][28] ),
    .A3(\soc/cpu/cpuregs/regs[7][28] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1600_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3124_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1600_ ),
    .Y(\soc/cpu/cpuregs/_1601_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3125_  (.A0(\soc/cpu/cpuregs/regs[0][28] ),
    .A1(\soc/cpu/cpuregs/regs[1][28] ),
    .A2(\soc/cpu/cpuregs/regs[4][28] ),
    .A3(\soc/cpu/cpuregs/regs[5][28] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1602_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3126_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1602_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1603_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3127_  (.A1(\soc/cpu/cpuregs/_1597_ ),
    .A2(\soc/cpu/cpuregs/_1599_ ),
    .B1(\soc/cpu/cpuregs/_1601_ ),
    .B2(\soc/cpu/cpuregs/_1603_ ),
    .Y(\soc/cpu/cpuregs/_1604_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3128_  (.A0(\soc/cpu/cpuregs/regs[24][28] ),
    .A1(\soc/cpu/cpuregs/regs[25][28] ),
    .A2(\soc/cpu/cpuregs/regs[28][28] ),
    .A3(\soc/cpu/cpuregs/regs[29][28] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1605_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3129_  (.A(net314),
    .B(\soc/cpu/cpuregs/_1605_ ),
    .Y(\soc/cpu/cpuregs/_1606_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3130_  (.A0(\soc/cpu/cpuregs/regs[26][28] ),
    .A1(\soc/cpu/cpuregs/regs[27][28] ),
    .A2(\soc/cpu/cpuregs/regs[30][28] ),
    .A3(\soc/cpu/cpuregs/regs[31][28] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1607_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3131_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1607_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1608_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3132_  (.A0(\soc/cpu/cpuregs/regs[10][28] ),
    .A1(\soc/cpu/cpuregs/regs[11][28] ),
    .A2(\soc/cpu/cpuregs/regs[14][28] ),
    .A3(\soc/cpu/cpuregs/regs[15][28] ),
    .S0(net322),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1609_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3133_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1609_ ),
    .Y(\soc/cpu/cpuregs/_1610_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3134_  (.A0(\soc/cpu/cpuregs/regs[8][28] ),
    .A1(\soc/cpu/cpuregs/regs[9][28] ),
    .A2(\soc/cpu/cpuregs/regs[12][28] ),
    .A3(\soc/cpu/cpuregs/regs[13][28] ),
    .S0(net320),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1611_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3135_  (.A1(net314),
    .A2(\soc/cpu/cpuregs/_1611_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1612_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3136_  (.A1(\soc/cpu/cpuregs/_1606_ ),
    .A2(\soc/cpu/cpuregs/_1608_ ),
    .B1(\soc/cpu/cpuregs/_1610_ ),
    .B2(\soc/cpu/cpuregs/_1612_ ),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1613_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3137_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1604_ ),
    .B1(\soc/cpu/cpuregs/_1613_ ),
    .X(\soc/cpu/cpuregs_rdata2[28] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3138_  (.A0(\soc/cpu/cpuregs/regs[16][29] ),
    .A1(\soc/cpu/cpuregs/regs[17][29] ),
    .A2(\soc/cpu/cpuregs/regs[20][29] ),
    .A3(\soc/cpu/cpuregs/regs[21][29] ),
    .S0(net326),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1614_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3139_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1614_ ),
    .Y(\soc/cpu/cpuregs/_1615_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3140_  (.A0(\soc/cpu/cpuregs/regs[18][29] ),
    .A1(\soc/cpu/cpuregs/regs[19][29] ),
    .A2(\soc/cpu/cpuregs/regs[22][29] ),
    .A3(\soc/cpu/cpuregs/regs[23][29] ),
    .S0(net326),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1616_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3141_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1616_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1617_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3142_  (.A0(\soc/cpu/cpuregs/regs[2][29] ),
    .A1(\soc/cpu/cpuregs/regs[3][29] ),
    .A2(\soc/cpu/cpuregs/regs[6][29] ),
    .A3(\soc/cpu/cpuregs/regs[7][29] ),
    .S0(net326),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1618_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3143_  (.A(net153),
    .B(\soc/cpu/cpuregs/_1618_ ),
    .Y(\soc/cpu/cpuregs/_1619_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3144_  (.A0(\soc/cpu/cpuregs/regs[0][29] ),
    .A1(\soc/cpu/cpuregs/regs[1][29] ),
    .A2(\soc/cpu/cpuregs/regs[4][29] ),
    .A3(\soc/cpu/cpuregs/regs[5][29] ),
    .S0(net324),
    .S1(\soc/cpu/cpuregs_raddr2[2] ),
    .X(\soc/cpu/cpuregs/_1620_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3145_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1620_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1621_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3146_  (.A1(\soc/cpu/cpuregs/_1615_ ),
    .A2(\soc/cpu/cpuregs/_1617_ ),
    .B1(\soc/cpu/cpuregs/_1619_ ),
    .B2(\soc/cpu/cpuregs/_1621_ ),
    .Y(\soc/cpu/cpuregs/_1622_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3147_  (.A0(\soc/cpu/cpuregs/regs[24][29] ),
    .A1(\soc/cpu/cpuregs/regs[25][29] ),
    .A2(\soc/cpu/cpuregs/regs[28][29] ),
    .A3(\soc/cpu/cpuregs/regs[29][29] ),
    .S0(net324),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1623_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3148_  (.A(net315),
    .B(\soc/cpu/cpuregs/_1623_ ),
    .Y(\soc/cpu/cpuregs/_1624_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3149_  (.A0(\soc/cpu/cpuregs/regs[26][29] ),
    .A1(\soc/cpu/cpuregs/regs[27][29] ),
    .A2(\soc/cpu/cpuregs/regs[30][29] ),
    .A3(\soc/cpu/cpuregs/regs[31][29] ),
    .S0(net324),
    .S1(net309),
    .X(\soc/cpu/cpuregs/_1625_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3150_  (.A1(net153),
    .A2(\soc/cpu/cpuregs/_1625_ ),
    .B1(net301),
    .Y(\soc/cpu/cpuregs/_1626_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3151_  (.A0(\soc/cpu/cpuregs/regs[10][29] ),
    .A1(\soc/cpu/cpuregs/regs[11][29] ),
    .A2(\soc/cpu/cpuregs/regs[14][29] ),
    .A3(\soc/cpu/cpuregs/regs[15][29] ),
    .S0(net324),
    .S1(net310),
    .X(\soc/cpu/cpuregs/_1627_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3152_  (.A0(\soc/cpu/cpuregs/regs[8][29] ),
    .A1(\soc/cpu/cpuregs/regs[9][29] ),
    .A2(\soc/cpu/cpuregs/regs[12][29] ),
    .A3(\soc/cpu/cpuregs/regs[13][29] ),
    .S0(net324),
    .S1(\soc/cpu/cpuregs_raddr2[2] ),
    .X(\soc/cpu/cpuregs/_1628_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3153_  (.A0(\soc/cpu/cpuregs/_1627_ ),
    .A1(\soc/cpu/cpuregs/_1628_ ),
    .S(net153),
    .Y(\soc/cpu/cpuregs/_1629_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3154_  (.A1(\soc/cpu/cpuregs/_1624_ ),
    .A2(\soc/cpu/cpuregs/_1626_ ),
    .B1(\soc/cpu/cpuregs/_1629_ ),
    .B2(net301),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1630_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3155_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1622_ ),
    .B1(\soc/cpu/cpuregs/_1630_ ),
    .X(\soc/cpu/cpuregs_rdata2[29] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3156_  (.A0(\soc/cpu/cpuregs/regs[26][30] ),
    .A1(\soc/cpu/cpuregs/regs[27][30] ),
    .A2(\soc/cpu/cpuregs/regs[30][30] ),
    .A3(\soc/cpu/cpuregs/regs[31][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1631_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3157_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1631_ ),
    .Y(\soc/cpu/cpuregs/_1632_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3158_  (.A0(\soc/cpu/cpuregs/regs[24][30] ),
    .A1(\soc/cpu/cpuregs/regs[25][30] ),
    .A2(\soc/cpu/cpuregs/regs[28][30] ),
    .A3(\soc/cpu/cpuregs/regs[29][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1633_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3159_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1633_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1634_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3160_  (.A0(\soc/cpu/cpuregs/regs[10][30] ),
    .A1(\soc/cpu/cpuregs/regs[11][30] ),
    .A2(\soc/cpu/cpuregs/regs[14][30] ),
    .A3(\soc/cpu/cpuregs/regs[15][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1635_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3161_  (.A0(\soc/cpu/cpuregs/regs[8][30] ),
    .A1(\soc/cpu/cpuregs/regs[9][30] ),
    .A2(\soc/cpu/cpuregs/regs[12][30] ),
    .A3(\soc/cpu/cpuregs/regs[13][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1636_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3162_  (.A0(\soc/cpu/cpuregs/_1635_ ),
    .A1(\soc/cpu/cpuregs/_1636_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1637_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3163_  (.A1(\soc/cpu/cpuregs/_1632_ ),
    .A2(\soc/cpu/cpuregs/_1634_ ),
    .B1(\soc/cpu/cpuregs/_1637_ ),
    .B2(net300),
    .Y(\soc/cpu/cpuregs/_1638_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3164_  (.A0(\soc/cpu/cpuregs/regs[2][30] ),
    .A1(\soc/cpu/cpuregs/regs[3][30] ),
    .A2(\soc/cpu/cpuregs/regs[6][30] ),
    .A3(\soc/cpu/cpuregs/regs[7][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1639_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3165_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1639_ ),
    .Y(\soc/cpu/cpuregs/_1640_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3166_  (.A0(\soc/cpu/cpuregs/regs[0][30] ),
    .A1(\soc/cpu/cpuregs/regs[1][30] ),
    .A2(\soc/cpu/cpuregs/regs[4][30] ),
    .A3(\soc/cpu/cpuregs/regs[5][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1641_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3167_  (.A1(net315),
    .A2(\soc/cpu/cpuregs/_1641_ ),
    .B1(\soc/cpu/cpuregs/_1059_ ),
    .Y(\soc/cpu/cpuregs/_1642_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3168_  (.A0(\soc/cpu/cpuregs/regs[18][30] ),
    .A1(\soc/cpu/cpuregs/regs[19][30] ),
    .A2(\soc/cpu/cpuregs/regs[22][30] ),
    .A3(\soc/cpu/cpuregs/regs[23][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1643_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3169_  (.A0(\soc/cpu/cpuregs/regs[16][30] ),
    .A1(\soc/cpu/cpuregs/regs[17][30] ),
    .A2(\soc/cpu/cpuregs/regs[20][30] ),
    .A3(\soc/cpu/cpuregs/regs[21][30] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1644_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3170_  (.A0(\soc/cpu/cpuregs/_1643_ ),
    .A1(\soc/cpu/cpuregs/_1644_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1645_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3171_  (.A1(\soc/cpu/cpuregs/_1640_ ),
    .A2(\soc/cpu/cpuregs/_1642_ ),
    .B1(\soc/cpu/cpuregs/_1645_ ),
    .B2(\soc/cpu/cpuregs/_1059_ ),
    .C1(\soc/cpu/cpuregs/_1025_ ),
    .Y(\soc/cpu/cpuregs/_1646_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3172_  (.A1(\soc/cpu/cpuregs/_1025_ ),
    .A2(\soc/cpu/cpuregs/_1638_ ),
    .B1(\soc/cpu/cpuregs/_1646_ ),
    .X(\soc/cpu/cpuregs_rdata2[30] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3173_  (.A0(\soc/cpu/cpuregs/regs[2][31] ),
    .A1(\soc/cpu/cpuregs/regs[3][31] ),
    .A2(\soc/cpu/cpuregs/regs[6][31] ),
    .A3(\soc/cpu/cpuregs/regs[7][31] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1647_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3174_  (.A(\soc/cpu/cpuregs/_1037_ ),
    .B(\soc/cpu/cpuregs/_1647_ ),
    .Y(\soc/cpu/cpuregs/_1648_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3175_  (.A0(\soc/cpu/cpuregs/regs[0][31] ),
    .A1(\soc/cpu/cpuregs/regs[1][31] ),
    .A2(\soc/cpu/cpuregs/regs[4][31] ),
    .A3(\soc/cpu/cpuregs/regs[5][31] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1649_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3176_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1649_ ),
    .Y(\soc/cpu/cpuregs/_1650_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3177_  (.A0(\soc/cpu/cpuregs/regs[16][31] ),
    .A1(\soc/cpu/cpuregs/regs[17][31] ),
    .A2(\soc/cpu/cpuregs/regs[20][31] ),
    .A3(\soc/cpu/cpuregs/regs[21][31] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1651_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3178_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1651_ ),
    .Y(\soc/cpu/cpuregs/_1652_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3179_  (.A0(\soc/cpu/cpuregs/regs[18][31] ),
    .A1(\soc/cpu/cpuregs/regs[19][31] ),
    .A2(\soc/cpu/cpuregs/regs[22][31] ),
    .A3(\soc/cpu/cpuregs/regs[23][31] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1653_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3180_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1653_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1654_ ));
 sky130_fd_sc_hd__o32ai_2 \soc/cpu/cpuregs/_3181_  (.A1(net300),
    .A2(\soc/cpu/cpuregs/_1648_ ),
    .A3(\soc/cpu/cpuregs/_1650_ ),
    .B1(\soc/cpu/cpuregs/_1652_ ),
    .B2(\soc/cpu/cpuregs/_1654_ ),
    .Y(\soc/cpu/cpuregs/_1655_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3182_  (.A0(\soc/cpu/cpuregs/regs[24][31] ),
    .A1(\soc/cpu/cpuregs/regs[25][31] ),
    .A2(\soc/cpu/cpuregs/regs[28][31] ),
    .A3(\soc/cpu/cpuregs/regs[29][31] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1656_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3183_  (.A(net313),
    .B(\soc/cpu/cpuregs/_1656_ ),
    .Y(\soc/cpu/cpuregs/_1657_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3184_  (.A0(\soc/cpu/cpuregs/regs[26][31] ),
    .A1(\soc/cpu/cpuregs/regs[27][31] ),
    .A2(\soc/cpu/cpuregs/regs[30][31] ),
    .A3(\soc/cpu/cpuregs/regs[31][31] ),
    .S0(net323),
    .S1(net311),
    .X(\soc/cpu/cpuregs/_1658_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_3185_  (.A1(\soc/cpu/cpuregs/_1037_ ),
    .A2(\soc/cpu/cpuregs/_1658_ ),
    .B1(net300),
    .Y(\soc/cpu/cpuregs/_1659_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3186_  (.A0(\soc/cpu/cpuregs/regs[10][31] ),
    .A1(\soc/cpu/cpuregs/regs[11][31] ),
    .A2(\soc/cpu/cpuregs/regs[14][31] ),
    .A3(\soc/cpu/cpuregs/regs[15][31] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1660_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3187_  (.A0(\soc/cpu/cpuregs/regs[8][31] ),
    .A1(\soc/cpu/cpuregs/regs[9][31] ),
    .A2(\soc/cpu/cpuregs/regs[12][31] ),
    .A3(\soc/cpu/cpuregs/regs[13][31] ),
    .S0(net325),
    .S1(net312),
    .X(\soc/cpu/cpuregs/_1661_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_3188_  (.A0(\soc/cpu/cpuregs/_1660_ ),
    .A1(\soc/cpu/cpuregs/_1661_ ),
    .S(\soc/cpu/cpuregs/_1037_ ),
    .Y(\soc/cpu/cpuregs/_1662_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3189_  (.A1(\soc/cpu/cpuregs/_1657_ ),
    .A2(\soc/cpu/cpuregs/_1659_ ),
    .B1(\soc/cpu/cpuregs/_1662_ ),
    .B2(net300),
    .C1(net303),
    .Y(\soc/cpu/cpuregs/_1663_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3190_  (.A1(net303),
    .A2(\soc/cpu/cpuregs/_1655_ ),
    .B1(\soc/cpu/cpuregs/_1663_ ),
    .X(\soc/cpu/cpuregs_rdata2[31] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3202_  (.A0(\soc/cpu/cpuregs/regs[16][0] ),
    .A1(\soc/cpu/cpuregs/regs[17][0] ),
    .A2(\soc/cpu/cpuregs/regs[20][0] ),
    .A3(\soc/cpu/cpuregs/regs[21][0] ),
    .S0(net351),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1675_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3203_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1675_ ),
    .Y(\soc/cpu/cpuregs/_1676_ ));
 sky130_fd_sc_hd__clkinv_16 \soc/cpu/cpuregs/_3204_  (.A(net342),
    .Y(\soc/cpu/cpuregs/_1677_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3210_  (.A0(\soc/cpu/cpuregs/regs[18][0] ),
    .A1(\soc/cpu/cpuregs/regs[19][0] ),
    .A2(\soc/cpu/cpuregs/regs[22][0] ),
    .A3(\soc/cpu/cpuregs/regs[23][0] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1683_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3213_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1683_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1686_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3219_  (.A0(\soc/cpu/cpuregs/regs[2][0] ),
    .A1(\soc/cpu/cpuregs/regs[3][0] ),
    .A2(\soc/cpu/cpuregs/regs[6][0] ),
    .A3(\soc/cpu/cpuregs/regs[7][0] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1692_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3220_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1692_ ),
    .Y(\soc/cpu/cpuregs/_1693_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3225_  (.A0(\soc/cpu/cpuregs/regs[0][0] ),
    .A1(\soc/cpu/cpuregs/regs[1][0] ),
    .A2(\soc/cpu/cpuregs/regs[4][0] ),
    .A3(\soc/cpu/cpuregs/regs[5][0] ),
    .S0(net351),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1698_ ));
 sky130_fd_sc_hd__clkinv_16 \soc/cpu/cpuregs/_3226_  (.A(net327),
    .Y(\soc/cpu/cpuregs/_1699_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3229_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_1698_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1702_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3230_  (.A1(\soc/cpu/cpuregs/_1676_ ),
    .A2(\soc/cpu/cpuregs/_1686_ ),
    .B1(\soc/cpu/cpuregs/_1693_ ),
    .B2(\soc/cpu/cpuregs/_1702_ ),
    .Y(\soc/cpu/cpuregs/_1703_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3235_  (.A0(\soc/cpu/cpuregs/regs[24][0] ),
    .A1(\soc/cpu/cpuregs/regs[25][0] ),
    .A2(\soc/cpu/cpuregs/regs[28][0] ),
    .A3(\soc/cpu/cpuregs/regs[29][0] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1708_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3236_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1708_ ),
    .Y(\soc/cpu/cpuregs/_1709_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3240_  (.A0(\soc/cpu/cpuregs/regs[26][0] ),
    .A1(\soc/cpu/cpuregs/regs[27][0] ),
    .A2(\soc/cpu/cpuregs/regs[30][0] ),
    .A3(\soc/cpu/cpuregs/regs[31][0] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1713_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_3242_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1713_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1715_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3248_  (.A0(\soc/cpu/cpuregs/regs[10][0] ),
    .A1(\soc/cpu/cpuregs/regs[11][0] ),
    .A2(\soc/cpu/cpuregs/regs[14][0] ),
    .A3(\soc/cpu/cpuregs/regs[15][0] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1721_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3249_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1721_ ),
    .Y(\soc/cpu/cpuregs/_1722_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3254_  (.A0(\soc/cpu/cpuregs/regs[8][0] ),
    .A1(\soc/cpu/cpuregs/regs[9][0] ),
    .A2(\soc/cpu/cpuregs/regs[12][0] ),
    .A3(\soc/cpu/cpuregs/regs[13][0] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1727_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3256_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_1727_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1729_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3259_  (.A1(\soc/cpu/cpuregs/_1709_ ),
    .A2(\soc/cpu/cpuregs/_1715_ ),
    .B1(\soc/cpu/cpuregs/_1722_ ),
    .B2(\soc/cpu/cpuregs/_1729_ ),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_1732_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3260_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_1703_ ),
    .B1(\soc/cpu/cpuregs/_1732_ ),
    .X(\soc/cpu/cpuregs_rdata1[0] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3262_  (.A0(\soc/cpu/cpuregs/regs[2][1] ),
    .A1(\soc/cpu/cpuregs/regs[3][1] ),
    .A2(\soc/cpu/cpuregs/regs[6][1] ),
    .A3(\soc/cpu/cpuregs/regs[7][1] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1734_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3264_  (.A0(\soc/cpu/cpuregs/regs[18][1] ),
    .A1(\soc/cpu/cpuregs/regs[19][1] ),
    .A2(\soc/cpu/cpuregs/regs[22][1] ),
    .A3(\soc/cpu/cpuregs/regs[23][1] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1736_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3266_  (.A0(\soc/cpu/cpuregs/regs[10][1] ),
    .A1(\soc/cpu/cpuregs/regs[11][1] ),
    .A2(\soc/cpu/cpuregs/regs[14][1] ),
    .A3(\soc/cpu/cpuregs/regs[15][1] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1738_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3269_  (.A0(\soc/cpu/cpuregs/regs[26][1] ),
    .A1(\soc/cpu/cpuregs/regs[27][1] ),
    .A2(\soc/cpu/cpuregs/regs[30][1] ),
    .A3(\soc/cpu/cpuregs/regs[31][1] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1741_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3270_  (.A0(\soc/cpu/cpuregs/_1734_ ),
    .A1(\soc/cpu/cpuregs/_1736_ ),
    .A2(\soc/cpu/cpuregs/_1738_ ),
    .A3(\soc/cpu/cpuregs/_1741_ ),
    .S0(net329),
    .S1(net331),
    .X(\soc/cpu/cpuregs/_1742_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3271_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1742_ ),
    .Y(\soc/cpu/cpuregs/_1743_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3273_  (.A0(\soc/cpu/cpuregs/regs[16][1] ),
    .A1(\soc/cpu/cpuregs/regs[17][1] ),
    .A2(\soc/cpu/cpuregs/regs[20][1] ),
    .A3(\soc/cpu/cpuregs/regs[21][1] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1745_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3274_  (.A0(\soc/cpu/cpuregs/regs[0][1] ),
    .A1(\soc/cpu/cpuregs/regs[1][1] ),
    .A2(\soc/cpu/cpuregs/regs[4][1] ),
    .A3(\soc/cpu/cpuregs/regs[5][1] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1746_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3275_  (.A0(\soc/cpu/cpuregs/regs[24][1] ),
    .A1(\soc/cpu/cpuregs/regs[25][1] ),
    .A2(\soc/cpu/cpuregs/regs[28][1] ),
    .A3(\soc/cpu/cpuregs/regs[29][1] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1747_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3276_  (.A0(\soc/cpu/cpuregs/regs[8][1] ),
    .A1(\soc/cpu/cpuregs/regs[9][1] ),
    .A2(\soc/cpu/cpuregs/regs[12][1] ),
    .A3(\soc/cpu/cpuregs/regs[13][1] ),
    .S0(net351),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1748_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3277_  (.A0(\soc/cpu/cpuregs/_1745_ ),
    .A1(\soc/cpu/cpuregs/_1746_ ),
    .A2(\soc/cpu/cpuregs/_1747_ ),
    .A3(\soc/cpu/cpuregs/_1748_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(net331),
    .X(\soc/cpu/cpuregs/_1749_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3278_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1749_ ),
    .Y(\soc/cpu/cpuregs/_1750_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/cpuregs/_3279_  (.A(\soc/cpu/cpuregs/_1743_ ),
    .B(\soc/cpu/cpuregs/_1750_ ),
    .Y(\soc/cpu/cpuregs_rdata1[1] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3280_  (.A0(\soc/cpu/cpuregs/regs[16][2] ),
    .A1(\soc/cpu/cpuregs/regs[17][2] ),
    .A2(\soc/cpu/cpuregs/regs[20][2] ),
    .A3(\soc/cpu/cpuregs/regs[21][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1751_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3281_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1751_ ),
    .Y(\soc/cpu/cpuregs/_1752_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3282_  (.A0(\soc/cpu/cpuregs/regs[18][2] ),
    .A1(\soc/cpu/cpuregs/regs[19][2] ),
    .A2(\soc/cpu/cpuregs/regs[22][2] ),
    .A3(\soc/cpu/cpuregs/regs[23][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1753_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3283_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1753_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1754_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3285_  (.A0(\soc/cpu/cpuregs/regs[2][2] ),
    .A1(\soc/cpu/cpuregs/regs[3][2] ),
    .A2(\soc/cpu/cpuregs/regs[6][2] ),
    .A3(\soc/cpu/cpuregs/regs[7][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1756_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3286_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1756_ ),
    .Y(\soc/cpu/cpuregs/_1757_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3287_  (.A0(\soc/cpu/cpuregs/regs[0][2] ),
    .A1(\soc/cpu/cpuregs/regs[1][2] ),
    .A2(\soc/cpu/cpuregs/regs[4][2] ),
    .A3(\soc/cpu/cpuregs/regs[5][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1758_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3288_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_1758_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1759_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3289_  (.A1(\soc/cpu/cpuregs/_1752_ ),
    .A2(\soc/cpu/cpuregs/_1754_ ),
    .B1(\soc/cpu/cpuregs/_1757_ ),
    .B2(\soc/cpu/cpuregs/_1759_ ),
    .Y(\soc/cpu/cpuregs/_1760_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3291_  (.A0(\soc/cpu/cpuregs/regs[24][2] ),
    .A1(\soc/cpu/cpuregs/regs[25][2] ),
    .A2(\soc/cpu/cpuregs/regs[28][2] ),
    .A3(\soc/cpu/cpuregs/regs[29][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1762_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3292_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1762_ ),
    .Y(\soc/cpu/cpuregs/_1763_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3293_  (.A0(\soc/cpu/cpuregs/regs[26][2] ),
    .A1(\soc/cpu/cpuregs/regs[27][2] ),
    .A2(\soc/cpu/cpuregs/regs[30][2] ),
    .A3(\soc/cpu/cpuregs/regs[31][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1764_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3294_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1764_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1765_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3297_  (.A0(\soc/cpu/cpuregs/regs[10][2] ),
    .A1(\soc/cpu/cpuregs/regs[11][2] ),
    .A2(\soc/cpu/cpuregs/regs[14][2] ),
    .A3(\soc/cpu/cpuregs/regs[15][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1768_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3300_  (.A0(\soc/cpu/cpuregs/regs[8][2] ),
    .A1(\soc/cpu/cpuregs/regs[9][2] ),
    .A2(\soc/cpu/cpuregs/regs[12][2] ),
    .A3(\soc/cpu/cpuregs/regs[13][2] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1771_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_3302_  (.A0(\soc/cpu/cpuregs/_1768_ ),
    .A1(\soc/cpu/cpuregs/_1771_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_1773_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3304_  (.A1(\soc/cpu/cpuregs/_1763_ ),
    .A2(\soc/cpu/cpuregs/_1765_ ),
    .B1(\soc/cpu/cpuregs/_1773_ ),
    .B2(net329),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_1775_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3305_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_1760_ ),
    .B1(\soc/cpu/cpuregs/_1775_ ),
    .X(\soc/cpu/cpuregs_rdata1[2] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3306_  (.A0(\soc/cpu/cpuregs/regs[16][3] ),
    .A1(\soc/cpu/cpuregs/regs[17][3] ),
    .A2(\soc/cpu/cpuregs/regs[20][3] ),
    .A3(\soc/cpu/cpuregs/regs[21][3] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1776_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3307_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1776_ ),
    .Y(\soc/cpu/cpuregs/_1777_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3308_  (.A0(\soc/cpu/cpuregs/regs[18][3] ),
    .A1(\soc/cpu/cpuregs/regs[19][3] ),
    .A2(\soc/cpu/cpuregs/regs[22][3] ),
    .A3(\soc/cpu/cpuregs/regs[23][3] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1778_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3309_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1778_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1779_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3310_  (.A0(\soc/cpu/cpuregs/regs[2][3] ),
    .A1(\soc/cpu/cpuregs/regs[3][3] ),
    .A2(\soc/cpu/cpuregs/regs[6][3] ),
    .A3(\soc/cpu/cpuregs/regs[7][3] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1780_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3311_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_1780_ ),
    .Y(\soc/cpu/cpuregs/_1781_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3313_  (.A0(\soc/cpu/cpuregs/regs[0][3] ),
    .A1(\soc/cpu/cpuregs/regs[1][3] ),
    .A2(\soc/cpu/cpuregs/regs[4][3] ),
    .A3(\soc/cpu/cpuregs/regs[5][3] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1783_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3314_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_1783_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1784_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3315_  (.A1(\soc/cpu/cpuregs/_1777_ ),
    .A2(\soc/cpu/cpuregs/_1779_ ),
    .B1(\soc/cpu/cpuregs/_1781_ ),
    .B2(\soc/cpu/cpuregs/_1784_ ),
    .Y(\soc/cpu/cpuregs/_1785_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3316_  (.A0(\soc/cpu/cpuregs/regs[24][3] ),
    .A1(\soc/cpu/cpuregs/regs[25][3] ),
    .A2(\soc/cpu/cpuregs/regs[28][3] ),
    .A3(\soc/cpu/cpuregs/regs[29][3] ),
    .S0(net349),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1786_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3317_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1786_ ),
    .Y(\soc/cpu/cpuregs/_1787_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3318_  (.A0(\soc/cpu/cpuregs/regs[26][3] ),
    .A1(\soc/cpu/cpuregs/regs[27][3] ),
    .A2(\soc/cpu/cpuregs/regs[30][3] ),
    .A3(\soc/cpu/cpuregs/regs[31][3] ),
    .S0(net349),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1788_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3319_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1788_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1789_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3320_  (.A0(\soc/cpu/cpuregs/regs[10][3] ),
    .A1(\soc/cpu/cpuregs/regs[11][3] ),
    .A2(\soc/cpu/cpuregs/regs[14][3] ),
    .A3(\soc/cpu/cpuregs/regs[15][3] ),
    .S0(net349),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_1790_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3322_  (.A0(\soc/cpu/cpuregs/regs[8][3] ),
    .A1(\soc/cpu/cpuregs/regs[9][3] ),
    .A2(\soc/cpu/cpuregs/regs[12][3] ),
    .A3(\soc/cpu/cpuregs/regs[13][3] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_1792_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3323_  (.A0(\soc/cpu/cpuregs/_1790_ ),
    .A1(\soc/cpu/cpuregs/_1792_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_1793_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3324_  (.A1(\soc/cpu/cpuregs/_1787_ ),
    .A2(\soc/cpu/cpuregs/_1789_ ),
    .B1(\soc/cpu/cpuregs/_1793_ ),
    .B2(net329),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_1794_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3325_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_1785_ ),
    .B1(\soc/cpu/cpuregs/_1794_ ),
    .X(\soc/cpu/cpuregs_rdata1[3] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3328_  (.A0(\soc/cpu/cpuregs/regs[2][4] ),
    .A1(\soc/cpu/cpuregs/regs[3][4] ),
    .A2(\soc/cpu/cpuregs/regs[6][4] ),
    .A3(\soc/cpu/cpuregs/regs[7][4] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_1797_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3329_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1797_ ),
    .Y(\soc/cpu/cpuregs/_1798_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3332_  (.A0(\soc/cpu/cpuregs/regs[0][4] ),
    .A1(\soc/cpu/cpuregs/regs[1][4] ),
    .A2(\soc/cpu/cpuregs/regs[4][4] ),
    .A3(\soc/cpu/cpuregs/regs[5][4] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_1801_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3333_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_1801_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1802_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3334_  (.A0(\soc/cpu/cpuregs/regs[16][4] ),
    .A1(\soc/cpu/cpuregs/regs[17][4] ),
    .A2(\soc/cpu/cpuregs/regs[20][4] ),
    .A3(\soc/cpu/cpuregs/regs[21][4] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_1803_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3335_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1803_ ),
    .Y(\soc/cpu/cpuregs/_1804_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3336_  (.A0(\soc/cpu/cpuregs/regs[18][4] ),
    .A1(\soc/cpu/cpuregs/regs[19][4] ),
    .A2(\soc/cpu/cpuregs/regs[22][4] ),
    .A3(\soc/cpu/cpuregs/regs[23][4] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1805_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3337_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1805_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_1806_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3338_  (.A1(\soc/cpu/cpuregs/_1798_ ),
    .A2(\soc/cpu/cpuregs/_1802_ ),
    .B1(\soc/cpu/cpuregs/_1804_ ),
    .B2(\soc/cpu/cpuregs/_1806_ ),
    .Y(\soc/cpu/cpuregs/_1807_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3339_  (.A0(\soc/cpu/cpuregs/regs[10][4] ),
    .A1(\soc/cpu/cpuregs/regs[11][4] ),
    .A2(\soc/cpu/cpuregs/regs[14][4] ),
    .A3(\soc/cpu/cpuregs/regs[15][4] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1808_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3340_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1808_ ),
    .Y(\soc/cpu/cpuregs/_1809_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3341_  (.A0(\soc/cpu/cpuregs/regs[8][4] ),
    .A1(\soc/cpu/cpuregs/regs[9][4] ),
    .A2(\soc/cpu/cpuregs/regs[12][4] ),
    .A3(\soc/cpu/cpuregs/regs[13][4] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1810_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3343_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_1810_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1812_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3344_  (.A0(\soc/cpu/cpuregs/regs[24][4] ),
    .A1(\soc/cpu/cpuregs/regs[25][4] ),
    .A2(\soc/cpu/cpuregs/regs[28][4] ),
    .A3(\soc/cpu/cpuregs/regs[29][4] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1813_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3345_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1813_ ),
    .Y(\soc/cpu/cpuregs/_1814_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3346_  (.A0(\soc/cpu/cpuregs/regs[26][4] ),
    .A1(\soc/cpu/cpuregs/regs[27][4] ),
    .A2(\soc/cpu/cpuregs/regs[30][4] ),
    .A3(\soc/cpu/cpuregs/regs[31][4] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1815_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_3348_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1815_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_1817_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3349_  (.A1(\soc/cpu/cpuregs/_1809_ ),
    .A2(\soc/cpu/cpuregs/_1812_ ),
    .B1(\soc/cpu/cpuregs/_1814_ ),
    .B2(\soc/cpu/cpuregs/_1817_ ),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_1818_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3350_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_1807_ ),
    .B1(\soc/cpu/cpuregs/_1818_ ),
    .X(\soc/cpu/cpuregs_rdata1[4] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3354_  (.A0(\soc/cpu/cpuregs/regs[2][5] ),
    .A1(\soc/cpu/cpuregs/regs[3][5] ),
    .A2(\soc/cpu/cpuregs/regs[6][5] ),
    .A3(\soc/cpu/cpuregs/regs[7][5] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_1822_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3355_  (.A0(\soc/cpu/cpuregs/regs[0][5] ),
    .A1(\soc/cpu/cpuregs/regs[1][5] ),
    .A2(\soc/cpu/cpuregs/regs[4][5] ),
    .A3(\soc/cpu/cpuregs/regs[5][5] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_1823_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3356_  (.A0(\soc/cpu/cpuregs/_1822_ ),
    .A1(\soc/cpu/cpuregs/_1823_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_1824_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3357_  (.A0(\soc/cpu/cpuregs/regs[16][5] ),
    .A1(\soc/cpu/cpuregs/regs[17][5] ),
    .A2(\soc/cpu/cpuregs/regs[20][5] ),
    .A3(\soc/cpu/cpuregs/regs[21][5] ),
    .S0(net352),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_1825_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3358_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1825_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1826_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3359_  (.A0(\soc/cpu/cpuregs/regs[18][5] ),
    .A1(\soc/cpu/cpuregs/regs[19][5] ),
    .A2(\soc/cpu/cpuregs/regs[22][5] ),
    .A3(\soc/cpu/cpuregs/regs[23][5] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1827_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_3360_  (.A(net342),
    .B(\soc/cpu/cpuregs/_1827_ ),
    .Y(\soc/cpu/cpuregs/_1828_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/cpuregs/_3361_  (.A1(\soc/cpu/cpuregs/_1699_ ),
    .A2(\soc/cpu/cpuregs/_1824_ ),
    .B1(\soc/cpu/cpuregs/_1826_ ),
    .B2(\soc/cpu/cpuregs/_1828_ ),
    .Y(\soc/cpu/cpuregs/_1829_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3363_  (.A0(\soc/cpu/cpuregs/regs[10][5] ),
    .A1(\soc/cpu/cpuregs/regs[11][5] ),
    .A2(\soc/cpu/cpuregs/regs[14][5] ),
    .A3(\soc/cpu/cpuregs/regs[15][5] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_1831_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3364_  (.A0(\soc/cpu/cpuregs/regs[8][5] ),
    .A1(\soc/cpu/cpuregs/regs[9][5] ),
    .A2(\soc/cpu/cpuregs/regs[12][5] ),
    .A3(\soc/cpu/cpuregs/regs[13][5] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1832_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3365_  (.A0(\soc/cpu/cpuregs/regs[26][5] ),
    .A1(\soc/cpu/cpuregs/regs[27][5] ),
    .A2(\soc/cpu/cpuregs/regs[30][5] ),
    .A3(\soc/cpu/cpuregs/regs[31][5] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1833_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3366_  (.A0(\soc/cpu/cpuregs/regs[24][5] ),
    .A1(\soc/cpu/cpuregs/regs[25][5] ),
    .A2(\soc/cpu/cpuregs/regs[28][5] ),
    .A3(\soc/cpu/cpuregs/regs[29][5] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1834_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3367_  (.A0(\soc/cpu/cpuregs/_1831_ ),
    .A1(\soc/cpu/cpuregs/_1832_ ),
    .A2(\soc/cpu/cpuregs/_1833_ ),
    .A3(\soc/cpu/cpuregs/_1834_ ),
    .S0(\soc/cpu/cpuregs/_1677_ ),
    .S1(net327),
    .X(\soc/cpu/cpuregs/_1835_ ));
 sky130_fd_sc_hd__mux2_4 \soc/cpu/cpuregs/_3368_  (.A0(\soc/cpu/cpuregs/_1829_ ),
    .A1(\soc/cpu/cpuregs/_1835_ ),
    .S(net332),
    .X(\soc/cpu/cpuregs_rdata1[5] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3369_  (.A0(\soc/cpu/cpuregs/regs[16][6] ),
    .A1(\soc/cpu/cpuregs/regs[17][6] ),
    .A2(\soc/cpu/cpuregs/regs[20][6] ),
    .A3(\soc/cpu/cpuregs/regs[21][6] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1836_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3370_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1836_ ),
    .Y(\soc/cpu/cpuregs/_1837_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3371_  (.A0(\soc/cpu/cpuregs/regs[18][6] ),
    .A1(\soc/cpu/cpuregs/regs[19][6] ),
    .A2(\soc/cpu/cpuregs/regs[22][6] ),
    .A3(\soc/cpu/cpuregs/regs[23][6] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1838_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3372_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1838_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1839_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3373_  (.A0(\soc/cpu/cpuregs/regs[2][6] ),
    .A1(\soc/cpu/cpuregs/regs[3][6] ),
    .A2(\soc/cpu/cpuregs/regs[6][6] ),
    .A3(\soc/cpu/cpuregs/regs[7][6] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1840_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3374_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1840_ ),
    .Y(\soc/cpu/cpuregs/_1841_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3376_  (.A0(\soc/cpu/cpuregs/regs[0][6] ),
    .A1(\soc/cpu/cpuregs/regs[1][6] ),
    .A2(\soc/cpu/cpuregs/regs[4][6] ),
    .A3(\soc/cpu/cpuregs/regs[5][6] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1843_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3377_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_1843_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1844_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3378_  (.A1(\soc/cpu/cpuregs/_1837_ ),
    .A2(\soc/cpu/cpuregs/_1839_ ),
    .B1(\soc/cpu/cpuregs/_1841_ ),
    .B2(\soc/cpu/cpuregs/_1844_ ),
    .Y(\soc/cpu/cpuregs/_1845_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3379_  (.A0(\soc/cpu/cpuregs/regs[24][6] ),
    .A1(\soc/cpu/cpuregs/regs[25][6] ),
    .A2(\soc/cpu/cpuregs/regs[28][6] ),
    .A3(\soc/cpu/cpuregs/regs[29][6] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1846_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3380_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1846_ ),
    .Y(\soc/cpu/cpuregs/_1847_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3382_  (.A0(\soc/cpu/cpuregs/regs[26][6] ),
    .A1(\soc/cpu/cpuregs/regs[27][6] ),
    .A2(\soc/cpu/cpuregs/regs[30][6] ),
    .A3(\soc/cpu/cpuregs/regs[31][6] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1849_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/cpu/cpuregs/_3383_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1849_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1850_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3384_  (.A0(\soc/cpu/cpuregs/regs[10][6] ),
    .A1(\soc/cpu/cpuregs/regs[11][6] ),
    .A2(\soc/cpu/cpuregs/regs[14][6] ),
    .A3(\soc/cpu/cpuregs/regs[15][6] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1851_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3385_  (.A0(\soc/cpu/cpuregs/regs[8][6] ),
    .A1(\soc/cpu/cpuregs/regs[9][6] ),
    .A2(\soc/cpu/cpuregs/regs[12][6] ),
    .A3(\soc/cpu/cpuregs/regs[13][6] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1852_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_3386_  (.A0(\soc/cpu/cpuregs/_1851_ ),
    .A1(\soc/cpu/cpuregs/_1852_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_1853_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3387_  (.A1(\soc/cpu/cpuregs/_1847_ ),
    .A2(\soc/cpu/cpuregs/_1850_ ),
    .B1(\soc/cpu/cpuregs/_1853_ ),
    .B2(net328),
    .C1(net330),
    .Y(\soc/cpu/cpuregs/_1854_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3388_  (.A1(net330),
    .A2(\soc/cpu/cpuregs/_1845_ ),
    .B1(\soc/cpu/cpuregs/_1854_ ),
    .X(\soc/cpu/cpuregs_rdata1[6] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3389_  (.A0(\soc/cpu/cpuregs/regs[16][7] ),
    .A1(\soc/cpu/cpuregs/regs[17][7] ),
    .A2(\soc/cpu/cpuregs/regs[20][7] ),
    .A3(\soc/cpu/cpuregs/regs[21][7] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1855_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3390_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1855_ ),
    .Y(\soc/cpu/cpuregs/_1856_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3391_  (.A0(\soc/cpu/cpuregs/regs[18][7] ),
    .A1(\soc/cpu/cpuregs/regs[19][7] ),
    .A2(\soc/cpu/cpuregs/regs[22][7] ),
    .A3(\soc/cpu/cpuregs/regs[23][7] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1857_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3392_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1857_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1858_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3393_  (.A0(\soc/cpu/cpuregs/regs[2][7] ),
    .A1(\soc/cpu/cpuregs/regs[3][7] ),
    .A2(\soc/cpu/cpuregs/regs[6][7] ),
    .A3(\soc/cpu/cpuregs/regs[7][7] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1859_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3394_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1859_ ),
    .Y(\soc/cpu/cpuregs/_1860_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3395_  (.A0(\soc/cpu/cpuregs/regs[0][7] ),
    .A1(\soc/cpu/cpuregs/regs[1][7] ),
    .A2(\soc/cpu/cpuregs/regs[4][7] ),
    .A3(\soc/cpu/cpuregs/regs[5][7] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1861_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3396_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_1861_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1862_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3397_  (.A1(\soc/cpu/cpuregs/_1856_ ),
    .A2(\soc/cpu/cpuregs/_1858_ ),
    .B1(\soc/cpu/cpuregs/_1860_ ),
    .B2(\soc/cpu/cpuregs/_1862_ ),
    .Y(\soc/cpu/cpuregs/_1863_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3398_  (.A0(\soc/cpu/cpuregs/regs[24][7] ),
    .A1(\soc/cpu/cpuregs/regs[25][7] ),
    .A2(\soc/cpu/cpuregs/regs[28][7] ),
    .A3(\soc/cpu/cpuregs/regs[29][7] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1864_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3399_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1864_ ),
    .Y(\soc/cpu/cpuregs/_1865_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3401_  (.A0(\soc/cpu/cpuregs/regs[26][7] ),
    .A1(\soc/cpu/cpuregs/regs[27][7] ),
    .A2(\soc/cpu/cpuregs/regs[30][7] ),
    .A3(\soc/cpu/cpuregs/regs[31][7] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1867_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3403_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1867_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1869_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3405_  (.A0(\soc/cpu/cpuregs/regs[10][7] ),
    .A1(\soc/cpu/cpuregs/regs[11][7] ),
    .A2(\soc/cpu/cpuregs/regs[14][7] ),
    .A3(\soc/cpu/cpuregs/regs[15][7] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1871_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3406_  (.A0(\soc/cpu/cpuregs/regs[8][7] ),
    .A1(\soc/cpu/cpuregs/regs[9][7] ),
    .A2(\soc/cpu/cpuregs/regs[12][7] ),
    .A3(\soc/cpu/cpuregs/regs[13][7] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1872_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_3407_  (.A0(\soc/cpu/cpuregs/_1871_ ),
    .A1(\soc/cpu/cpuregs/_1872_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_1873_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3408_  (.A1(\soc/cpu/cpuregs/_1865_ ),
    .A2(\soc/cpu/cpuregs/_1869_ ),
    .B1(\soc/cpu/cpuregs/_1873_ ),
    .B2(net328),
    .C1(net330),
    .Y(\soc/cpu/cpuregs/_1874_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3409_  (.A1(net330),
    .A2(\soc/cpu/cpuregs/_1863_ ),
    .B1(\soc/cpu/cpuregs/_1874_ ),
    .X(\soc/cpu/cpuregs_rdata1[7] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3410_  (.A0(\soc/cpu/cpuregs/regs[2][8] ),
    .A1(\soc/cpu/cpuregs/regs[3][8] ),
    .A2(\soc/cpu/cpuregs/regs[6][8] ),
    .A3(\soc/cpu/cpuregs/regs[7][8] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1875_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3411_  (.A0(\soc/cpu/cpuregs/regs[18][8] ),
    .A1(\soc/cpu/cpuregs/regs[19][8] ),
    .A2(\soc/cpu/cpuregs/regs[22][8] ),
    .A3(\soc/cpu/cpuregs/regs[23][8] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1876_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3412_  (.A0(\soc/cpu/cpuregs/regs[10][8] ),
    .A1(\soc/cpu/cpuregs/regs[11][8] ),
    .A2(\soc/cpu/cpuregs/regs[14][8] ),
    .A3(\soc/cpu/cpuregs/regs[15][8] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1877_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3413_  (.A0(\soc/cpu/cpuregs/regs[26][8] ),
    .A1(\soc/cpu/cpuregs/regs[27][8] ),
    .A2(\soc/cpu/cpuregs/regs[30][8] ),
    .A3(\soc/cpu/cpuregs/regs[31][8] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1878_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3414_  (.A0(\soc/cpu/cpuregs/_1875_ ),
    .A1(\soc/cpu/cpuregs/_1876_ ),
    .A2(\soc/cpu/cpuregs/_1877_ ),
    .A3(\soc/cpu/cpuregs/_1878_ ),
    .S0(net328),
    .S1(net330),
    .X(\soc/cpu/cpuregs/_1879_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3415_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1879_ ),
    .Y(\soc/cpu/cpuregs/_1880_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3416_  (.A0(\soc/cpu/cpuregs/regs[16][8] ),
    .A1(\soc/cpu/cpuregs/regs[17][8] ),
    .A2(\soc/cpu/cpuregs/regs[20][8] ),
    .A3(\soc/cpu/cpuregs/regs[21][8] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1881_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3417_  (.A0(\soc/cpu/cpuregs/regs[0][8] ),
    .A1(\soc/cpu/cpuregs/regs[1][8] ),
    .A2(\soc/cpu/cpuregs/regs[4][8] ),
    .A3(\soc/cpu/cpuregs/regs[5][8] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1882_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3418_  (.A0(\soc/cpu/cpuregs/regs[24][8] ),
    .A1(\soc/cpu/cpuregs/regs[25][8] ),
    .A2(\soc/cpu/cpuregs/regs[28][8] ),
    .A3(\soc/cpu/cpuregs/regs[29][8] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1883_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3419_  (.A0(\soc/cpu/cpuregs/regs[8][8] ),
    .A1(\soc/cpu/cpuregs/regs[9][8] ),
    .A2(\soc/cpu/cpuregs/regs[12][8] ),
    .A3(\soc/cpu/cpuregs/regs[13][8] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1884_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3420_  (.A0(\soc/cpu/cpuregs/_1881_ ),
    .A1(\soc/cpu/cpuregs/_1882_ ),
    .A2(\soc/cpu/cpuregs/_1883_ ),
    .A3(\soc/cpu/cpuregs/_1884_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(net330),
    .X(\soc/cpu/cpuregs/_1885_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3421_  (.A(net343),
    .B(\soc/cpu/cpuregs/_1885_ ),
    .Y(\soc/cpu/cpuregs/_1886_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/cpuregs/_3422_  (.A(\soc/cpu/cpuregs/_1880_ ),
    .B(\soc/cpu/cpuregs/_1886_ ),
    .Y(\soc/cpu/cpuregs_rdata1[8] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3423_  (.A0(\soc/cpu/cpuregs/regs[2][9] ),
    .A1(\soc/cpu/cpuregs/regs[3][9] ),
    .A2(\soc/cpu/cpuregs/regs[6][9] ),
    .A3(\soc/cpu/cpuregs/regs[7][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1887_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3424_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_1887_ ),
    .Y(\soc/cpu/cpuregs/_1888_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3425_  (.A0(\soc/cpu/cpuregs/regs[0][9] ),
    .A1(\soc/cpu/cpuregs/regs[1][9] ),
    .A2(\soc/cpu/cpuregs/regs[4][9] ),
    .A3(\soc/cpu/cpuregs/regs[5][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1889_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3426_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_1889_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1890_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3428_  (.A0(\soc/cpu/cpuregs/regs[16][9] ),
    .A1(\soc/cpu/cpuregs/regs[17][9] ),
    .A2(\soc/cpu/cpuregs/regs[20][9] ),
    .A3(\soc/cpu/cpuregs/regs[21][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1892_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3429_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1892_ ),
    .Y(\soc/cpu/cpuregs/_1893_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3430_  (.A0(\soc/cpu/cpuregs/regs[18][9] ),
    .A1(\soc/cpu/cpuregs/regs[19][9] ),
    .A2(\soc/cpu/cpuregs/regs[22][9] ),
    .A3(\soc/cpu/cpuregs/regs[23][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1894_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3431_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1894_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1895_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3432_  (.A1(\soc/cpu/cpuregs/_1888_ ),
    .A2(\soc/cpu/cpuregs/_1890_ ),
    .B1(\soc/cpu/cpuregs/_1893_ ),
    .B2(\soc/cpu/cpuregs/_1895_ ),
    .Y(\soc/cpu/cpuregs/_1896_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3434_  (.A0(\soc/cpu/cpuregs/regs[10][9] ),
    .A1(\soc/cpu/cpuregs/regs[11][9] ),
    .A2(\soc/cpu/cpuregs/regs[14][9] ),
    .A3(\soc/cpu/cpuregs/regs[15][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1898_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3435_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_1898_ ),
    .Y(\soc/cpu/cpuregs/_1899_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3437_  (.A0(\soc/cpu/cpuregs/regs[8][9] ),
    .A1(\soc/cpu/cpuregs/regs[9][9] ),
    .A2(\soc/cpu/cpuregs/regs[12][9] ),
    .A3(\soc/cpu/cpuregs/regs[13][9] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1901_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3438_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_1901_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1902_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3439_  (.A0(\soc/cpu/cpuregs/regs[24][9] ),
    .A1(\soc/cpu/cpuregs/regs[25][9] ),
    .A2(\soc/cpu/cpuregs/regs[28][9] ),
    .A3(\soc/cpu/cpuregs/regs[29][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1903_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3440_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1903_ ),
    .Y(\soc/cpu/cpuregs/_1904_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3441_  (.A0(\soc/cpu/cpuregs/regs[26][9] ),
    .A1(\soc/cpu/cpuregs/regs[27][9] ),
    .A2(\soc/cpu/cpuregs/regs[30][9] ),
    .A3(\soc/cpu/cpuregs/regs[31][9] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1905_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3442_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1905_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1906_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3443_  (.A1(\soc/cpu/cpuregs/_1899_ ),
    .A2(\soc/cpu/cpuregs/_1902_ ),
    .B1(\soc/cpu/cpuregs/_1904_ ),
    .B2(\soc/cpu/cpuregs/_1906_ ),
    .C1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_1907_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/cpuregs/_3444_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_1896_ ),
    .B1(\soc/cpu/cpuregs/_1907_ ),
    .X(\soc/cpu/cpuregs_rdata1[9] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3445_  (.A0(\soc/cpu/cpuregs/regs[16][10] ),
    .A1(\soc/cpu/cpuregs/regs[17][10] ),
    .A2(\soc/cpu/cpuregs/regs[20][10] ),
    .A3(\soc/cpu/cpuregs/regs[21][10] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1908_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3446_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1908_ ),
    .Y(\soc/cpu/cpuregs/_1909_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3447_  (.A0(\soc/cpu/cpuregs/regs[18][10] ),
    .A1(\soc/cpu/cpuregs/regs[19][10] ),
    .A2(\soc/cpu/cpuregs/regs[22][10] ),
    .A3(\soc/cpu/cpuregs/regs[23][10] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1910_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3448_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1910_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1911_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3450_  (.A0(\soc/cpu/cpuregs/regs[2][10] ),
    .A1(\soc/cpu/cpuregs/regs[3][10] ),
    .A2(\soc/cpu/cpuregs/regs[6][10] ),
    .A3(\soc/cpu/cpuregs/regs[7][10] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1913_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3451_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_1913_ ),
    .Y(\soc/cpu/cpuregs/_1914_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3452_  (.A0(\soc/cpu/cpuregs/regs[0][10] ),
    .A1(\soc/cpu/cpuregs/regs[1][10] ),
    .A2(\soc/cpu/cpuregs/regs[4][10] ),
    .A3(\soc/cpu/cpuregs/regs[5][10] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1915_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3453_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_1915_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1916_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3454_  (.A1(\soc/cpu/cpuregs/_1909_ ),
    .A2(\soc/cpu/cpuregs/_1911_ ),
    .B1(\soc/cpu/cpuregs/_1914_ ),
    .B2(\soc/cpu/cpuregs/_1916_ ),
    .Y(\soc/cpu/cpuregs/_1917_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3456_  (.A0(\soc/cpu/cpuregs/regs[24][10] ),
    .A1(\soc/cpu/cpuregs/regs[25][10] ),
    .A2(\soc/cpu/cpuregs/regs[28][10] ),
    .A3(\soc/cpu/cpuregs/regs[29][10] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_1919_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3457_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1919_ ),
    .Y(\soc/cpu/cpuregs/_1920_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3458_  (.A0(\soc/cpu/cpuregs/regs[26][10] ),
    .A1(\soc/cpu/cpuregs/regs[27][10] ),
    .A2(\soc/cpu/cpuregs/regs[30][10] ),
    .A3(\soc/cpu/cpuregs/regs[31][10] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1921_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3459_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1921_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1922_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3460_  (.A0(\soc/cpu/cpuregs/regs[10][10] ),
    .A1(\soc/cpu/cpuregs/regs[11][10] ),
    .A2(\soc/cpu/cpuregs/regs[14][10] ),
    .A3(\soc/cpu/cpuregs/regs[15][10] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1923_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3461_  (.A0(\soc/cpu/cpuregs/regs[8][10] ),
    .A1(\soc/cpu/cpuregs/regs[9][10] ),
    .A2(\soc/cpu/cpuregs/regs[12][10] ),
    .A3(\soc/cpu/cpuregs/regs[13][10] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1924_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3462_  (.A0(\soc/cpu/cpuregs/_1923_ ),
    .A1(\soc/cpu/cpuregs/_1924_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_1925_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3464_  (.A1(\soc/cpu/cpuregs/_1920_ ),
    .A2(\soc/cpu/cpuregs/_1922_ ),
    .B1(\soc/cpu/cpuregs/_1925_ ),
    .B2(net328),
    .C1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_1927_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3465_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_1917_ ),
    .B1(\soc/cpu/cpuregs/_1927_ ),
    .X(\soc/cpu/cpuregs_rdata1[10] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3467_  (.A0(\soc/cpu/cpuregs/regs[2][11] ),
    .A1(\soc/cpu/cpuregs/regs[3][11] ),
    .A2(\soc/cpu/cpuregs/regs[6][11] ),
    .A3(\soc/cpu/cpuregs/regs[7][11] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1929_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3468_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1929_ ),
    .Y(\soc/cpu/cpuregs/_1930_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3469_  (.A0(\soc/cpu/cpuregs/regs[0][11] ),
    .A1(\soc/cpu/cpuregs/regs[1][11] ),
    .A2(\soc/cpu/cpuregs/regs[4][11] ),
    .A3(\soc/cpu/cpuregs/regs[5][11] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1931_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3470_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_1931_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1932_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3471_  (.A0(\soc/cpu/cpuregs/regs[16][11] ),
    .A1(\soc/cpu/cpuregs/regs[17][11] ),
    .A2(\soc/cpu/cpuregs/regs[20][11] ),
    .A3(\soc/cpu/cpuregs/regs[21][11] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1933_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3472_  (.A(net343),
    .B(\soc/cpu/cpuregs/_1933_ ),
    .Y(\soc/cpu/cpuregs/_1934_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3474_  (.A0(\soc/cpu/cpuregs/regs[18][11] ),
    .A1(\soc/cpu/cpuregs/regs[19][11] ),
    .A2(\soc/cpu/cpuregs/regs[22][11] ),
    .A3(\soc/cpu/cpuregs/regs[23][11] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1936_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3475_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1936_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_1937_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3476_  (.A1(\soc/cpu/cpuregs/_1930_ ),
    .A2(\soc/cpu/cpuregs/_1932_ ),
    .B1(\soc/cpu/cpuregs/_1934_ ),
    .B2(\soc/cpu/cpuregs/_1937_ ),
    .Y(\soc/cpu/cpuregs/_1938_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3477_  (.A0(\soc/cpu/cpuregs/regs[10][11] ),
    .A1(\soc/cpu/cpuregs/regs[11][11] ),
    .A2(\soc/cpu/cpuregs/regs[14][11] ),
    .A3(\soc/cpu/cpuregs/regs[15][11] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1939_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3478_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1939_ ),
    .Y(\soc/cpu/cpuregs/_1940_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3479_  (.A0(\soc/cpu/cpuregs/regs[8][11] ),
    .A1(\soc/cpu/cpuregs/regs[9][11] ),
    .A2(\soc/cpu/cpuregs/regs[12][11] ),
    .A3(\soc/cpu/cpuregs/regs[13][11] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1941_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3480_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_1941_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1942_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3481_  (.A0(\soc/cpu/cpuregs/regs[24][11] ),
    .A1(\soc/cpu/cpuregs/regs[25][11] ),
    .A2(\soc/cpu/cpuregs/regs[28][11] ),
    .A3(\soc/cpu/cpuregs/regs[29][11] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1943_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3482_  (.A(net343),
    .B(\soc/cpu/cpuregs/_1943_ ),
    .Y(\soc/cpu/cpuregs/_1944_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3483_  (.A0(\soc/cpu/cpuregs/regs[26][11] ),
    .A1(\soc/cpu/cpuregs/regs[27][11] ),
    .A2(\soc/cpu/cpuregs/regs[30][11] ),
    .A3(\soc/cpu/cpuregs/regs[31][11] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_1945_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3484_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1945_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_1946_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3485_  (.A1(\soc/cpu/cpuregs/_1940_ ),
    .A2(\soc/cpu/cpuregs/_1942_ ),
    .B1(\soc/cpu/cpuregs/_1944_ ),
    .B2(\soc/cpu/cpuregs/_1946_ ),
    .C1(net332),
    .Y(\soc/cpu/cpuregs/_1947_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3486_  (.A1(net332),
    .A2(\soc/cpu/cpuregs/_1938_ ),
    .B1(\soc/cpu/cpuregs/_1947_ ),
    .X(\soc/cpu/cpuregs_rdata1[11] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3487_  (.A0(\soc/cpu/cpuregs/regs[2][12] ),
    .A1(\soc/cpu/cpuregs/regs[3][12] ),
    .A2(\soc/cpu/cpuregs/regs[6][12] ),
    .A3(\soc/cpu/cpuregs/regs[7][12] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1948_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3488_  (.A0(\soc/cpu/cpuregs/regs[18][12] ),
    .A1(\soc/cpu/cpuregs/regs[19][12] ),
    .A2(\soc/cpu/cpuregs/regs[22][12] ),
    .A3(\soc/cpu/cpuregs/regs[23][12] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1949_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3489_  (.A0(\soc/cpu/cpuregs/regs[10][12] ),
    .A1(\soc/cpu/cpuregs/regs[11][12] ),
    .A2(\soc/cpu/cpuregs/regs[14][12] ),
    .A3(\soc/cpu/cpuregs/regs[15][12] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1950_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3490_  (.A0(\soc/cpu/cpuregs/regs[26][12] ),
    .A1(\soc/cpu/cpuregs/regs[27][12] ),
    .A2(\soc/cpu/cpuregs/regs[30][12] ),
    .A3(\soc/cpu/cpuregs/regs[31][12] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1951_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3491_  (.A0(\soc/cpu/cpuregs/_1948_ ),
    .A1(\soc/cpu/cpuregs/_1949_ ),
    .A2(\soc/cpu/cpuregs/_1950_ ),
    .A3(\soc/cpu/cpuregs/_1951_ ),
    .S0(net328),
    .S1(\soc/cpu/cpuregs_raddr1[3] ),
    .X(\soc/cpu/cpuregs/_1952_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3492_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_1952_ ),
    .Y(\soc/cpu/cpuregs/_1953_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3493_  (.A0(\soc/cpu/cpuregs/regs[16][12] ),
    .A1(\soc/cpu/cpuregs/regs[17][12] ),
    .A2(\soc/cpu/cpuregs/regs[20][12] ),
    .A3(\soc/cpu/cpuregs/regs[21][12] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1954_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3494_  (.A0(\soc/cpu/cpuregs/regs[0][12] ),
    .A1(\soc/cpu/cpuregs/regs[1][12] ),
    .A2(\soc/cpu/cpuregs/regs[4][12] ),
    .A3(\soc/cpu/cpuregs/regs[5][12] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_1955_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3495_  (.A0(\soc/cpu/cpuregs/regs[24][12] ),
    .A1(\soc/cpu/cpuregs/regs[25][12] ),
    .A2(\soc/cpu/cpuregs/regs[28][12] ),
    .A3(\soc/cpu/cpuregs/regs[29][12] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1956_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3496_  (.A0(\soc/cpu/cpuregs/regs[8][12] ),
    .A1(\soc/cpu/cpuregs/regs[9][12] ),
    .A2(\soc/cpu/cpuregs/regs[12][12] ),
    .A3(\soc/cpu/cpuregs/regs[13][12] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1957_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3497_  (.A0(\soc/cpu/cpuregs/_1954_ ),
    .A1(\soc/cpu/cpuregs/_1955_ ),
    .A2(\soc/cpu/cpuregs/_1956_ ),
    .A3(\soc/cpu/cpuregs/_1957_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(\soc/cpu/cpuregs_raddr1[3] ),
    .X(\soc/cpu/cpuregs/_1958_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3498_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1958_ ),
    .Y(\soc/cpu/cpuregs/_1959_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_3499_  (.A(\soc/cpu/cpuregs/_1953_ ),
    .B(\soc/cpu/cpuregs/_1959_ ),
    .Y(\soc/cpu/cpuregs_rdata1[12] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3500_  (.A0(\soc/cpu/cpuregs/regs[16][13] ),
    .A1(\soc/cpu/cpuregs/regs[17][13] ),
    .A2(\soc/cpu/cpuregs/regs[20][13] ),
    .A3(\soc/cpu/cpuregs/regs[21][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1960_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3501_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1960_ ),
    .Y(\soc/cpu/cpuregs/_1961_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3504_  (.A0(\soc/cpu/cpuregs/regs[18][13] ),
    .A1(\soc/cpu/cpuregs/regs[19][13] ),
    .A2(\soc/cpu/cpuregs/regs[22][13] ),
    .A3(\soc/cpu/cpuregs/regs[23][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1964_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3505_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_1964_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1965_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3506_  (.A0(\soc/cpu/cpuregs/regs[2][13] ),
    .A1(\soc/cpu/cpuregs/regs[3][13] ),
    .A2(\soc/cpu/cpuregs/regs[6][13] ),
    .A3(\soc/cpu/cpuregs/regs[7][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1966_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3507_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_1966_ ),
    .Y(\soc/cpu/cpuregs/_1967_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3508_  (.A0(\soc/cpu/cpuregs/regs[0][13] ),
    .A1(\soc/cpu/cpuregs/regs[1][13] ),
    .A2(\soc/cpu/cpuregs/regs[4][13] ),
    .A3(\soc/cpu/cpuregs/regs[5][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1968_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3509_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_1968_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1969_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3510_  (.A1(\soc/cpu/cpuregs/_1961_ ),
    .A2(\soc/cpu/cpuregs/_1965_ ),
    .B1(\soc/cpu/cpuregs/_1967_ ),
    .B2(\soc/cpu/cpuregs/_1969_ ),
    .Y(\soc/cpu/cpuregs/_1970_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3511_  (.A0(\soc/cpu/cpuregs/regs[24][13] ),
    .A1(\soc/cpu/cpuregs/regs[25][13] ),
    .A2(\soc/cpu/cpuregs/regs[28][13] ),
    .A3(\soc/cpu/cpuregs/regs[29][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1971_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3512_  (.A(net341),
    .B(\soc/cpu/cpuregs/_1971_ ),
    .Y(\soc/cpu/cpuregs/_1972_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3513_  (.A0(\soc/cpu/cpuregs/regs[26][13] ),
    .A1(\soc/cpu/cpuregs/regs[27][13] ),
    .A2(\soc/cpu/cpuregs/regs[30][13] ),
    .A3(\soc/cpu/cpuregs/regs[31][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1973_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3514_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1973_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_1974_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3515_  (.A0(\soc/cpu/cpuregs/regs[10][13] ),
    .A1(\soc/cpu/cpuregs/regs[11][13] ),
    .A2(\soc/cpu/cpuregs/regs[14][13] ),
    .A3(\soc/cpu/cpuregs/regs[15][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1975_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3516_  (.A0(\soc/cpu/cpuregs/regs[8][13] ),
    .A1(\soc/cpu/cpuregs/regs[9][13] ),
    .A2(\soc/cpu/cpuregs/regs[12][13] ),
    .A3(\soc/cpu/cpuregs/regs[13][13] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_1976_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_3518_  (.A0(\soc/cpu/cpuregs/_1975_ ),
    .A1(\soc/cpu/cpuregs/_1976_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_1978_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3519_  (.A1(\soc/cpu/cpuregs/_1972_ ),
    .A2(\soc/cpu/cpuregs/_1974_ ),
    .B1(\soc/cpu/cpuregs/_1978_ ),
    .B2(net328),
    .C1(net330),
    .Y(\soc/cpu/cpuregs/_1979_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3520_  (.A1(net330),
    .A2(\soc/cpu/cpuregs/_1970_ ),
    .B1(\soc/cpu/cpuregs/_1979_ ),
    .X(\soc/cpu/cpuregs_rdata1[13] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3522_  (.A0(\soc/cpu/cpuregs/regs[16][14] ),
    .A1(\soc/cpu/cpuregs/regs[17][14] ),
    .A2(\soc/cpu/cpuregs/regs[20][14] ),
    .A3(\soc/cpu/cpuregs/regs[21][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1981_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3523_  (.A(net343),
    .B(\soc/cpu/cpuregs/_1981_ ),
    .Y(\soc/cpu/cpuregs/_1982_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3524_  (.A0(\soc/cpu/cpuregs/regs[18][14] ),
    .A1(\soc/cpu/cpuregs/regs[19][14] ),
    .A2(\soc/cpu/cpuregs/regs[22][14] ),
    .A3(\soc/cpu/cpuregs/regs[23][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1983_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3526_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1983_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1985_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3527_  (.A0(\soc/cpu/cpuregs/regs[2][14] ),
    .A1(\soc/cpu/cpuregs/regs[3][14] ),
    .A2(\soc/cpu/cpuregs/regs[6][14] ),
    .A3(\soc/cpu/cpuregs/regs[7][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1986_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3528_  (.A(net152),
    .B(\soc/cpu/cpuregs/_1986_ ),
    .Y(\soc/cpu/cpuregs/_1987_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3529_  (.A0(\soc/cpu/cpuregs/regs[0][14] ),
    .A1(\soc/cpu/cpuregs/regs[1][14] ),
    .A2(\soc/cpu/cpuregs/regs[4][14] ),
    .A3(\soc/cpu/cpuregs/regs[5][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1988_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3530_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_1988_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_1989_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3531_  (.A1(\soc/cpu/cpuregs/_1982_ ),
    .A2(\soc/cpu/cpuregs/_1985_ ),
    .B1(\soc/cpu/cpuregs/_1987_ ),
    .B2(\soc/cpu/cpuregs/_1989_ ),
    .Y(\soc/cpu/cpuregs/_1990_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3532_  (.A0(\soc/cpu/cpuregs/regs[24][14] ),
    .A1(\soc/cpu/cpuregs/regs[25][14] ),
    .A2(\soc/cpu/cpuregs/regs[28][14] ),
    .A3(\soc/cpu/cpuregs/regs[29][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1991_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3533_  (.A(net343),
    .B(\soc/cpu/cpuregs/_1991_ ),
    .Y(\soc/cpu/cpuregs/_1992_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3534_  (.A0(\soc/cpu/cpuregs/regs[26][14] ),
    .A1(\soc/cpu/cpuregs/regs[27][14] ),
    .A2(\soc/cpu/cpuregs/regs[30][14] ),
    .A3(\soc/cpu/cpuregs/regs[31][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1993_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3535_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_1993_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_1994_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3536_  (.A0(\soc/cpu/cpuregs/regs[10][14] ),
    .A1(\soc/cpu/cpuregs/regs[11][14] ),
    .A2(\soc/cpu/cpuregs/regs[14][14] ),
    .A3(\soc/cpu/cpuregs/regs[15][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1995_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3537_  (.A0(\soc/cpu/cpuregs/regs[8][14] ),
    .A1(\soc/cpu/cpuregs/regs[9][14] ),
    .A2(\soc/cpu/cpuregs/regs[12][14] ),
    .A3(\soc/cpu/cpuregs/regs[13][14] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_1996_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_3538_  (.A0(\soc/cpu/cpuregs/_1995_ ),
    .A1(\soc/cpu/cpuregs/_1996_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_1997_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3539_  (.A1(\soc/cpu/cpuregs/_1992_ ),
    .A2(\soc/cpu/cpuregs/_1994_ ),
    .B1(\soc/cpu/cpuregs/_1997_ ),
    .B2(net329),
    .C1(net332),
    .Y(\soc/cpu/cpuregs/_1998_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3540_  (.A1(net332),
    .A2(\soc/cpu/cpuregs/_1990_ ),
    .B1(\soc/cpu/cpuregs/_1998_ ),
    .X(\soc/cpu/cpuregs_rdata1[14] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3541_  (.A0(\soc/cpu/cpuregs/regs[18][15] ),
    .A1(\soc/cpu/cpuregs/regs[19][15] ),
    .A2(\soc/cpu/cpuregs/regs[22][15] ),
    .A3(\soc/cpu/cpuregs/regs[23][15] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_1999_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3542_  (.A0(\soc/cpu/cpuregs/regs[26][15] ),
    .A1(\soc/cpu/cpuregs/regs[27][15] ),
    .A2(\soc/cpu/cpuregs/regs[30][15] ),
    .A3(\soc/cpu/cpuregs/regs[31][15] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2000_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3543_  (.A0(\soc/cpu/cpuregs/_1999_ ),
    .A1(\soc/cpu/cpuregs/_2000_ ),
    .S(net330),
    .X(\soc/cpu/cpuregs/_2001_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3544_  (.A(\soc/cpu/cpuregs/_1699_ ),
    .B(\soc/cpu/cpuregs/_2001_ ),
    .Y(\soc/cpu/cpuregs/_2002_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3545_  (.A0(\soc/cpu/cpuregs/regs[10][15] ),
    .A1(\soc/cpu/cpuregs/regs[11][15] ),
    .A2(\soc/cpu/cpuregs/regs[14][15] ),
    .A3(\soc/cpu/cpuregs/regs[15][15] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2003_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/cpuregs/_3546_  (.A(\soc/cpu/cpuregs/regs[2][15] ),
    .SLEEP(net334),
    .X(\soc/cpu/cpuregs/_2004_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/cpuregs/_3547_  (.A1(\soc/cpu/cpuregs/regs[6][15] ),
    .A2(net334),
    .B1(\soc/cpu/cpuregs/_2004_ ),
    .C1(net345),
    .X(\soc/cpu/cpuregs/_2005_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3548_  (.A0(\soc/cpu/cpuregs/regs[3][15] ),
    .A1(\soc/cpu/cpuregs/regs[7][15] ),
    .S(net334),
    .Y(\soc/cpu/cpuregs/_2006_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3549_  (.A1(net345),
    .A2(\soc/cpu/cpuregs/_2006_ ),
    .B1(net330),
    .Y(\soc/cpu/cpuregs/_2007_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/cpu/cpuregs/_3550_  (.A1(net330),
    .A2(\soc/cpu/cpuregs/_2003_ ),
    .B1(\soc/cpu/cpuregs/_2005_ ),
    .B2(\soc/cpu/cpuregs/_2007_ ),
    .C1(net328),
    .Y(\soc/cpu/cpuregs/_2008_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3551_  (.A0(\soc/cpu/cpuregs/regs[16][15] ),
    .A1(\soc/cpu/cpuregs/regs[17][15] ),
    .A2(\soc/cpu/cpuregs/regs[20][15] ),
    .A3(\soc/cpu/cpuregs/regs[21][15] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2009_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3552_  (.A0(\soc/cpu/cpuregs/regs[0][15] ),
    .A1(\soc/cpu/cpuregs/regs[1][15] ),
    .A2(\soc/cpu/cpuregs/regs[4][15] ),
    .A3(\soc/cpu/cpuregs/regs[5][15] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2010_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3553_  (.A0(\soc/cpu/cpuregs/regs[24][15] ),
    .A1(\soc/cpu/cpuregs/regs[25][15] ),
    .A2(\soc/cpu/cpuregs/regs[28][15] ),
    .A3(\soc/cpu/cpuregs/regs[29][15] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2011_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3554_  (.A0(\soc/cpu/cpuregs/regs[8][15] ),
    .A1(\soc/cpu/cpuregs/regs[9][15] ),
    .A2(\soc/cpu/cpuregs/regs[12][15] ),
    .A3(\soc/cpu/cpuregs/regs[13][15] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2012_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3555_  (.A0(\soc/cpu/cpuregs/_2009_ ),
    .A1(\soc/cpu/cpuregs/_2010_ ),
    .A2(\soc/cpu/cpuregs/_2011_ ),
    .A3(\soc/cpu/cpuregs/_2012_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(net330),
    .X(\soc/cpu/cpuregs/_2013_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_3556_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2013_ ),
    .Y(\soc/cpu/cpuregs/_2014_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/cpu/cpuregs/_3557_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2002_ ),
    .A3(\soc/cpu/cpuregs/_2008_ ),
    .B1(\soc/cpu/cpuregs/_2014_ ),
    .Y(\soc/cpu/cpuregs_rdata1[15] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3558_  (.A0(\soc/cpu/cpuregs/regs[2][16] ),
    .A1(\soc/cpu/cpuregs/regs[3][16] ),
    .A2(\soc/cpu/cpuregs/regs[6][16] ),
    .A3(\soc/cpu/cpuregs/regs[7][16] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2015_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3559_  (.A0(\soc/cpu/cpuregs/regs[18][16] ),
    .A1(\soc/cpu/cpuregs/regs[19][16] ),
    .A2(\soc/cpu/cpuregs/regs[22][16] ),
    .A3(\soc/cpu/cpuregs/regs[23][16] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2016_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3560_  (.A0(\soc/cpu/cpuregs/regs[10][16] ),
    .A1(\soc/cpu/cpuregs/regs[11][16] ),
    .A2(\soc/cpu/cpuregs/regs[14][16] ),
    .A3(\soc/cpu/cpuregs/regs[15][16] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2017_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3561_  (.A0(\soc/cpu/cpuregs/regs[26][16] ),
    .A1(\soc/cpu/cpuregs/regs[27][16] ),
    .A2(\soc/cpu/cpuregs/regs[30][16] ),
    .A3(\soc/cpu/cpuregs/regs[31][16] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2018_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3562_  (.A0(\soc/cpu/cpuregs/_2015_ ),
    .A1(\soc/cpu/cpuregs/_2016_ ),
    .A2(\soc/cpu/cpuregs/_2017_ ),
    .A3(\soc/cpu/cpuregs/_2018_ ),
    .S0(net328),
    .S1(\soc/cpu/cpuregs_raddr1[3] ),
    .X(\soc/cpu/cpuregs/_2019_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3563_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2019_ ),
    .Y(\soc/cpu/cpuregs/_2020_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3564_  (.A0(\soc/cpu/cpuregs/regs[16][16] ),
    .A1(\soc/cpu/cpuregs/regs[17][16] ),
    .A2(\soc/cpu/cpuregs/regs[20][16] ),
    .A3(\soc/cpu/cpuregs/regs[21][16] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2021_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3565_  (.A0(\soc/cpu/cpuregs/regs[0][16] ),
    .A1(\soc/cpu/cpuregs/regs[1][16] ),
    .A2(\soc/cpu/cpuregs/regs[4][16] ),
    .A3(\soc/cpu/cpuregs/regs[5][16] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2022_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3566_  (.A0(\soc/cpu/cpuregs/regs[24][16] ),
    .A1(\soc/cpu/cpuregs/regs[25][16] ),
    .A2(\soc/cpu/cpuregs/regs[28][16] ),
    .A3(\soc/cpu/cpuregs/regs[29][16] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2023_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3567_  (.A0(\soc/cpu/cpuregs/regs[8][16] ),
    .A1(\soc/cpu/cpuregs/regs[9][16] ),
    .A2(\soc/cpu/cpuregs/regs[12][16] ),
    .A3(\soc/cpu/cpuregs/regs[13][16] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2024_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3568_  (.A0(\soc/cpu/cpuregs/_2021_ ),
    .A1(\soc/cpu/cpuregs/_2022_ ),
    .A2(\soc/cpu/cpuregs/_2023_ ),
    .A3(\soc/cpu/cpuregs/_2024_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(\soc/cpu/cpuregs_raddr1[3] ),
    .X(\soc/cpu/cpuregs/_2025_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3569_  (.A(net341),
    .B(\soc/cpu/cpuregs/_2025_ ),
    .Y(\soc/cpu/cpuregs/_2026_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_3570_  (.A(\soc/cpu/cpuregs/_2020_ ),
    .B(\soc/cpu/cpuregs/_2026_ ),
    .Y(\soc/cpu/cpuregs_rdata1[16] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3571_  (.A0(\soc/cpu/cpuregs/regs[2][17] ),
    .A1(\soc/cpu/cpuregs/regs[3][17] ),
    .A2(\soc/cpu/cpuregs/regs[6][17] ),
    .A3(\soc/cpu/cpuregs/regs[7][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2027_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3572_  (.A0(\soc/cpu/cpuregs/regs[18][17] ),
    .A1(\soc/cpu/cpuregs/regs[19][17] ),
    .A2(\soc/cpu/cpuregs/regs[22][17] ),
    .A3(\soc/cpu/cpuregs/regs[23][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2028_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3573_  (.A0(\soc/cpu/cpuregs/regs[10][17] ),
    .A1(\soc/cpu/cpuregs/regs[11][17] ),
    .A2(\soc/cpu/cpuregs/regs[14][17] ),
    .A3(\soc/cpu/cpuregs/regs[15][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2029_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3574_  (.A0(\soc/cpu/cpuregs/regs[26][17] ),
    .A1(\soc/cpu/cpuregs/regs[27][17] ),
    .A2(\soc/cpu/cpuregs/regs[30][17] ),
    .A3(\soc/cpu/cpuregs/regs[31][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2030_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3575_  (.A0(\soc/cpu/cpuregs/_2027_ ),
    .A1(\soc/cpu/cpuregs/_2028_ ),
    .A2(\soc/cpu/cpuregs/_2029_ ),
    .A3(\soc/cpu/cpuregs/_2030_ ),
    .S0(net327),
    .S1(net330),
    .X(\soc/cpu/cpuregs/_2031_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_3576_  (.A(net152),
    .B(\soc/cpu/cpuregs/_2031_ ),
    .Y(\soc/cpu/cpuregs/_2032_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3577_  (.A0(\soc/cpu/cpuregs/regs[16][17] ),
    .A1(\soc/cpu/cpuregs/regs[17][17] ),
    .A2(\soc/cpu/cpuregs/regs[20][17] ),
    .A3(\soc/cpu/cpuregs/regs[21][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2033_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3578_  (.A0(\soc/cpu/cpuregs/regs[0][17] ),
    .A1(\soc/cpu/cpuregs/regs[1][17] ),
    .A2(\soc/cpu/cpuregs/regs[4][17] ),
    .A3(\soc/cpu/cpuregs/regs[5][17] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2034_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3579_  (.A0(\soc/cpu/cpuregs/regs[24][17] ),
    .A1(\soc/cpu/cpuregs/regs[25][17] ),
    .A2(\soc/cpu/cpuregs/regs[28][17] ),
    .A3(\soc/cpu/cpuregs/regs[29][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2035_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3580_  (.A0(\soc/cpu/cpuregs/regs[8][17] ),
    .A1(\soc/cpu/cpuregs/regs[9][17] ),
    .A2(\soc/cpu/cpuregs/regs[12][17] ),
    .A3(\soc/cpu/cpuregs/regs[13][17] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2036_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3581_  (.A0(\soc/cpu/cpuregs/_2033_ ),
    .A1(\soc/cpu/cpuregs/_2034_ ),
    .A2(\soc/cpu/cpuregs/_2035_ ),
    .A3(\soc/cpu/cpuregs/_2036_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(net330),
    .X(\soc/cpu/cpuregs/_2037_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_3582_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2037_ ),
    .Y(\soc/cpu/cpuregs/_2038_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_3583_  (.A(\soc/cpu/cpuregs/_2032_ ),
    .B(\soc/cpu/cpuregs/_2038_ ),
    .Y(\soc/cpu/cpuregs_rdata1[17] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3584_  (.A0(\soc/cpu/cpuregs/regs[16][18] ),
    .A1(\soc/cpu/cpuregs/regs[17][18] ),
    .A2(\soc/cpu/cpuregs/regs[20][18] ),
    .A3(\soc/cpu/cpuregs/regs[21][18] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2039_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3585_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2039_ ),
    .Y(\soc/cpu/cpuregs/_2040_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3586_  (.A0(\soc/cpu/cpuregs/regs[18][18] ),
    .A1(\soc/cpu/cpuregs/regs[19][18] ),
    .A2(\soc/cpu/cpuregs/regs[22][18] ),
    .A3(\soc/cpu/cpuregs/regs[23][18] ),
    .S0(net353),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2041_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3587_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2041_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2042_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3589_  (.A0(\soc/cpu/cpuregs/regs[2][18] ),
    .A1(\soc/cpu/cpuregs/regs[3][18] ),
    .A2(\soc/cpu/cpuregs/regs[6][18] ),
    .A3(\soc/cpu/cpuregs/regs[7][18] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2044_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3590_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2044_ ),
    .Y(\soc/cpu/cpuregs/_2045_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3591_  (.A0(\soc/cpu/cpuregs/regs[0][18] ),
    .A1(\soc/cpu/cpuregs/regs[1][18] ),
    .A2(\soc/cpu/cpuregs/regs[4][18] ),
    .A3(\soc/cpu/cpuregs/regs[5][18] ),
    .S0(net353),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2046_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3592_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_2046_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2047_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3593_  (.A1(\soc/cpu/cpuregs/_2040_ ),
    .A2(\soc/cpu/cpuregs/_2042_ ),
    .B1(\soc/cpu/cpuregs/_2045_ ),
    .B2(\soc/cpu/cpuregs/_2047_ ),
    .Y(\soc/cpu/cpuregs/_2048_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3594_  (.A0(\soc/cpu/cpuregs/regs[24][18] ),
    .A1(\soc/cpu/cpuregs/regs[25][18] ),
    .A2(\soc/cpu/cpuregs/regs[28][18] ),
    .A3(\soc/cpu/cpuregs/regs[29][18] ),
    .S0(net352),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2049_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3595_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2049_ ),
    .Y(\soc/cpu/cpuregs/_2050_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3596_  (.A0(\soc/cpu/cpuregs/regs[26][18] ),
    .A1(\soc/cpu/cpuregs/regs[27][18] ),
    .A2(\soc/cpu/cpuregs/regs[30][18] ),
    .A3(\soc/cpu/cpuregs/regs[31][18] ),
    .S0(net352),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2051_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3597_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2051_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_2052_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3598_  (.A0(\soc/cpu/cpuregs/regs[10][18] ),
    .A1(\soc/cpu/cpuregs/regs[11][18] ),
    .A2(\soc/cpu/cpuregs/regs[14][18] ),
    .A3(\soc/cpu/cpuregs/regs[15][18] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2053_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3599_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2053_ ),
    .Y(\soc/cpu/cpuregs/_2054_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3600_  (.A0(\soc/cpu/cpuregs/regs[8][18] ),
    .A1(\soc/cpu/cpuregs/regs[9][18] ),
    .A2(\soc/cpu/cpuregs/regs[12][18] ),
    .A3(\soc/cpu/cpuregs/regs[13][18] ),
    .S0(net352),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2055_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3601_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_2055_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2056_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3602_  (.A1(\soc/cpu/cpuregs/_2050_ ),
    .A2(\soc/cpu/cpuregs/_2052_ ),
    .B1(\soc/cpu/cpuregs/_2054_ ),
    .B2(\soc/cpu/cpuregs/_2056_ ),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_2057_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3603_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_2048_ ),
    .B1(\soc/cpu/cpuregs/_2057_ ),
    .X(\soc/cpu/cpuregs_rdata1[18] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3604_  (.A0(\soc/cpu/cpuregs/regs[16][19] ),
    .A1(\soc/cpu/cpuregs/regs[17][19] ),
    .A2(\soc/cpu/cpuregs/regs[20][19] ),
    .A3(\soc/cpu/cpuregs/regs[21][19] ),
    .S0(net353),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2058_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3605_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2058_ ),
    .Y(\soc/cpu/cpuregs/_2059_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3606_  (.A0(\soc/cpu/cpuregs/regs[18][19] ),
    .A1(\soc/cpu/cpuregs/regs[19][19] ),
    .A2(\soc/cpu/cpuregs/regs[22][19] ),
    .A3(\soc/cpu/cpuregs/regs[23][19] ),
    .S0(net353),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2060_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3607_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2060_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2061_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3608_  (.A0(\soc/cpu/cpuregs/regs[2][19] ),
    .A1(\soc/cpu/cpuregs/regs[3][19] ),
    .A2(\soc/cpu/cpuregs/regs[6][19] ),
    .A3(\soc/cpu/cpuregs/regs[7][19] ),
    .S0(net353),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2062_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3609_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2062_ ),
    .Y(\soc/cpu/cpuregs/_2063_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3611_  (.A0(\soc/cpu/cpuregs/regs[0][19] ),
    .A1(\soc/cpu/cpuregs/regs[1][19] ),
    .A2(\soc/cpu/cpuregs/regs[4][19] ),
    .A3(\soc/cpu/cpuregs/regs[5][19] ),
    .S0(net353),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2065_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3612_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_2065_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2066_ ));
 sky130_fd_sc_hd__o22ai_4 \soc/cpu/cpuregs/_3613_  (.A1(\soc/cpu/cpuregs/_2059_ ),
    .A2(\soc/cpu/cpuregs/_2061_ ),
    .B1(\soc/cpu/cpuregs/_2063_ ),
    .B2(\soc/cpu/cpuregs/_2066_ ),
    .Y(\soc/cpu/cpuregs/_2067_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3614_  (.A0(\soc/cpu/cpuregs/regs[24][19] ),
    .A1(\soc/cpu/cpuregs/regs[25][19] ),
    .A2(\soc/cpu/cpuregs/regs[28][19] ),
    .A3(\soc/cpu/cpuregs/regs[29][19] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2068_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3615_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2068_ ),
    .Y(\soc/cpu/cpuregs/_2069_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3616_  (.A0(\soc/cpu/cpuregs/regs[26][19] ),
    .A1(\soc/cpu/cpuregs/regs[27][19] ),
    .A2(\soc/cpu/cpuregs/regs[30][19] ),
    .A3(\soc/cpu/cpuregs/regs[31][19] ),
    .S0(net352),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2070_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3617_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2070_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_2071_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3618_  (.A0(\soc/cpu/cpuregs/regs[10][19] ),
    .A1(\soc/cpu/cpuregs/regs[11][19] ),
    .A2(\soc/cpu/cpuregs/regs[14][19] ),
    .A3(\soc/cpu/cpuregs/regs[15][19] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2072_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3619_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2072_ ),
    .Y(\soc/cpu/cpuregs/_2073_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3620_  (.A0(\soc/cpu/cpuregs/regs[8][19] ),
    .A1(\soc/cpu/cpuregs/regs[9][19] ),
    .A2(\soc/cpu/cpuregs/regs[12][19] ),
    .A3(\soc/cpu/cpuregs/regs[13][19] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2074_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3621_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2074_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2075_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3622_  (.A1(\soc/cpu/cpuregs/_2069_ ),
    .A2(\soc/cpu/cpuregs/_2071_ ),
    .B1(\soc/cpu/cpuregs/_2073_ ),
    .B2(\soc/cpu/cpuregs/_2075_ ),
    .C1(net332),
    .Y(\soc/cpu/cpuregs/_2076_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3623_  (.A1(net332),
    .A2(\soc/cpu/cpuregs/_2067_ ),
    .B1(\soc/cpu/cpuregs/_2076_ ),
    .X(\soc/cpu/cpuregs_rdata1[19] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3624_  (.A0(\soc/cpu/cpuregs/regs[2][20] ),
    .A1(\soc/cpu/cpuregs/regs[3][20] ),
    .A2(\soc/cpu/cpuregs/regs[6][20] ),
    .A3(\soc/cpu/cpuregs/regs[7][20] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2077_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3625_  (.A0(\soc/cpu/cpuregs/regs[18][20] ),
    .A1(\soc/cpu/cpuregs/regs[19][20] ),
    .A2(\soc/cpu/cpuregs/regs[22][20] ),
    .A3(\soc/cpu/cpuregs/regs[23][20] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2078_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3626_  (.A0(\soc/cpu/cpuregs/regs[10][20] ),
    .A1(\soc/cpu/cpuregs/regs[11][20] ),
    .A2(\soc/cpu/cpuregs/regs[14][20] ),
    .A3(\soc/cpu/cpuregs/regs[15][20] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2079_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3627_  (.A0(\soc/cpu/cpuregs/regs[26][20] ),
    .A1(\soc/cpu/cpuregs/regs[27][20] ),
    .A2(\soc/cpu/cpuregs/regs[30][20] ),
    .A3(\soc/cpu/cpuregs/regs[31][20] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2080_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3628_  (.A0(\soc/cpu/cpuregs/_2077_ ),
    .A1(\soc/cpu/cpuregs/_2078_ ),
    .A2(\soc/cpu/cpuregs/_2079_ ),
    .A3(\soc/cpu/cpuregs/_2080_ ),
    .S0(net329),
    .S1(net332),
    .X(\soc/cpu/cpuregs/_2081_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3629_  (.A(net152),
    .B(\soc/cpu/cpuregs/_2081_ ),
    .Y(\soc/cpu/cpuregs/_2082_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3630_  (.A0(\soc/cpu/cpuregs/regs[16][20] ),
    .A1(\soc/cpu/cpuregs/regs[17][20] ),
    .A2(\soc/cpu/cpuregs/regs[20][20] ),
    .A3(\soc/cpu/cpuregs/regs[21][20] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2083_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3631_  (.A0(\soc/cpu/cpuregs/regs[0][20] ),
    .A1(\soc/cpu/cpuregs/regs[1][20] ),
    .A2(\soc/cpu/cpuregs/regs[4][20] ),
    .A3(\soc/cpu/cpuregs/regs[5][20] ),
    .S0(net350),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2084_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3632_  (.A0(\soc/cpu/cpuregs/regs[24][20] ),
    .A1(\soc/cpu/cpuregs/regs[25][20] ),
    .A2(\soc/cpu/cpuregs/regs[28][20] ),
    .A3(\soc/cpu/cpuregs/regs[29][20] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2085_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3633_  (.A0(\soc/cpu/cpuregs/regs[8][20] ),
    .A1(\soc/cpu/cpuregs/regs[9][20] ),
    .A2(\soc/cpu/cpuregs/regs[12][20] ),
    .A3(\soc/cpu/cpuregs/regs[13][20] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2086_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3634_  (.A0(\soc/cpu/cpuregs/_2083_ ),
    .A1(\soc/cpu/cpuregs/_2084_ ),
    .A2(\soc/cpu/cpuregs/_2085_ ),
    .A3(\soc/cpu/cpuregs/_2086_ ),
    .S0(\soc/cpu/cpuregs/_1699_ ),
    .S1(net332),
    .X(\soc/cpu/cpuregs/_2087_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3635_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2087_ ),
    .Y(\soc/cpu/cpuregs/_2088_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/cpuregs/_3636_  (.A(\soc/cpu/cpuregs/_2082_ ),
    .B(\soc/cpu/cpuregs/_2088_ ),
    .Y(\soc/cpu/cpuregs_rdata1[20] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3637_  (.A0(\soc/cpu/cpuregs/regs[2][21] ),
    .A1(\soc/cpu/cpuregs/regs[3][21] ),
    .A2(\soc/cpu/cpuregs/regs[6][21] ),
    .A3(\soc/cpu/cpuregs/regs[7][21] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2089_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3639_  (.A0(\soc/cpu/cpuregs/regs[0][21] ),
    .A1(\soc/cpu/cpuregs/regs[1][21] ),
    .A2(\soc/cpu/cpuregs/regs[4][21] ),
    .A3(\soc/cpu/cpuregs/regs[5][21] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2091_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3640_  (.A0(\soc/cpu/cpuregs/_2089_ ),
    .A1(\soc/cpu/cpuregs/_2091_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2092_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3641_  (.A0(\soc/cpu/cpuregs/regs[16][21] ),
    .A1(\soc/cpu/cpuregs/regs[17][21] ),
    .A2(\soc/cpu/cpuregs/regs[20][21] ),
    .A3(\soc/cpu/cpuregs/regs[21][21] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2093_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3642_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2093_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2094_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3643_  (.A0(\soc/cpu/cpuregs/regs[18][21] ),
    .A1(\soc/cpu/cpuregs/regs[19][21] ),
    .A2(\soc/cpu/cpuregs/regs[22][21] ),
    .A3(\soc/cpu/cpuregs/regs[23][21] ),
    .S0(net353),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2095_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_3644_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2095_ ),
    .Y(\soc/cpu/cpuregs/_2096_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/cpu/cpuregs/_3645_  (.A1(\soc/cpu/cpuregs/_1699_ ),
    .A2(\soc/cpu/cpuregs/_2092_ ),
    .B1(\soc/cpu/cpuregs/_2094_ ),
    .B2(\soc/cpu/cpuregs/_2096_ ),
    .Y(\soc/cpu/cpuregs/_2097_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3646_  (.A0(\soc/cpu/cpuregs/regs[10][21] ),
    .A1(\soc/cpu/cpuregs/regs[11][21] ),
    .A2(\soc/cpu/cpuregs/regs[14][21] ),
    .A3(\soc/cpu/cpuregs/regs[15][21] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2098_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3647_  (.A0(\soc/cpu/cpuregs/regs[8][21] ),
    .A1(\soc/cpu/cpuregs/regs[9][21] ),
    .A2(\soc/cpu/cpuregs/regs[12][21] ),
    .A3(\soc/cpu/cpuregs/regs[13][21] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2099_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3648_  (.A0(\soc/cpu/cpuregs/_2098_ ),
    .A1(\soc/cpu/cpuregs/_2099_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2100_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3649_  (.A0(\soc/cpu/cpuregs/regs[26][21] ),
    .A1(\soc/cpu/cpuregs/regs[27][21] ),
    .A2(\soc/cpu/cpuregs/regs[30][21] ),
    .A3(\soc/cpu/cpuregs/regs[31][21] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2101_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3650_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2101_ ),
    .Y(\soc/cpu/cpuregs/_2102_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3651_  (.A0(\soc/cpu/cpuregs/regs[24][21] ),
    .A1(\soc/cpu/cpuregs/regs[25][21] ),
    .A2(\soc/cpu/cpuregs/regs[28][21] ),
    .A3(\soc/cpu/cpuregs/regs[29][21] ),
    .S0(net351),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2103_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3652_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_2103_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_2104_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3653_  (.A1(net327),
    .A2(\soc/cpu/cpuregs/_2100_ ),
    .B1(\soc/cpu/cpuregs/_2102_ ),
    .B2(\soc/cpu/cpuregs/_2104_ ),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_2105_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3654_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_2097_ ),
    .B1(\soc/cpu/cpuregs/_2105_ ),
    .X(\soc/cpu/cpuregs_rdata1[21] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3655_  (.A0(\soc/cpu/cpuregs/regs[16][22] ),
    .A1(\soc/cpu/cpuregs/regs[17][22] ),
    .A2(\soc/cpu/cpuregs/regs[20][22] ),
    .A3(\soc/cpu/cpuregs/regs[21][22] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2106_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3656_  (.A(net341),
    .B(\soc/cpu/cpuregs/_2106_ ),
    .Y(\soc/cpu/cpuregs/_2107_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3657_  (.A0(\soc/cpu/cpuregs/regs[18][22] ),
    .A1(\soc/cpu/cpuregs/regs[19][22] ),
    .A2(\soc/cpu/cpuregs/regs[22][22] ),
    .A3(\soc/cpu/cpuregs/regs[23][22] ),
    .S0(net347),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2108_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3658_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2108_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2109_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3659_  (.A0(\soc/cpu/cpuregs/regs[2][22] ),
    .A1(\soc/cpu/cpuregs/regs[3][22] ),
    .A2(\soc/cpu/cpuregs/regs[6][22] ),
    .A3(\soc/cpu/cpuregs/regs[7][22] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2110_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3660_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2110_ ),
    .Y(\soc/cpu/cpuregs/_2111_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3661_  (.A0(\soc/cpu/cpuregs/regs[0][22] ),
    .A1(\soc/cpu/cpuregs/regs[1][22] ),
    .A2(\soc/cpu/cpuregs/regs[4][22] ),
    .A3(\soc/cpu/cpuregs/regs[5][22] ),
    .S0(net347),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2112_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3662_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_2112_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2113_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3663_  (.A1(\soc/cpu/cpuregs/_2107_ ),
    .A2(\soc/cpu/cpuregs/_2109_ ),
    .B1(\soc/cpu/cpuregs/_2111_ ),
    .B2(\soc/cpu/cpuregs/_2113_ ),
    .Y(\soc/cpu/cpuregs/_2114_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3664_  (.A0(\soc/cpu/cpuregs/regs[24][22] ),
    .A1(\soc/cpu/cpuregs/regs[25][22] ),
    .A2(\soc/cpu/cpuregs/regs[28][22] ),
    .A3(\soc/cpu/cpuregs/regs[29][22] ),
    .S0(net347),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2115_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3665_  (.A(net341),
    .B(\soc/cpu/cpuregs/_2115_ ),
    .Y(\soc/cpu/cpuregs/_2116_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3666_  (.A0(\soc/cpu/cpuregs/regs[26][22] ),
    .A1(\soc/cpu/cpuregs/regs[27][22] ),
    .A2(\soc/cpu/cpuregs/regs[30][22] ),
    .A3(\soc/cpu/cpuregs/regs[31][22] ),
    .S0(net346),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2117_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3667_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2117_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2118_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3668_  (.A0(\soc/cpu/cpuregs/regs[10][22] ),
    .A1(\soc/cpu/cpuregs/regs[11][22] ),
    .A2(\soc/cpu/cpuregs/regs[14][22] ),
    .A3(\soc/cpu/cpuregs/regs[15][22] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2119_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3669_  (.A0(\soc/cpu/cpuregs/regs[8][22] ),
    .A1(\soc/cpu/cpuregs/regs[9][22] ),
    .A2(\soc/cpu/cpuregs/regs[12][22] ),
    .A3(\soc/cpu/cpuregs/regs[13][22] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2120_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_3670_  (.A0(\soc/cpu/cpuregs/_2119_ ),
    .A1(\soc/cpu/cpuregs/_2120_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2121_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3671_  (.A1(\soc/cpu/cpuregs/_2116_ ),
    .A2(\soc/cpu/cpuregs/_2118_ ),
    .B1(\soc/cpu/cpuregs/_2121_ ),
    .B2(net328),
    .C1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_2122_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/cpuregs/_3672_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_2114_ ),
    .B1(\soc/cpu/cpuregs/_2122_ ),
    .X(\soc/cpu/cpuregs_rdata1[22] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3673_  (.A0(\soc/cpu/cpuregs/regs[16][23] ),
    .A1(\soc/cpu/cpuregs/regs[17][23] ),
    .A2(\soc/cpu/cpuregs/regs[20][23] ),
    .A3(\soc/cpu/cpuregs/regs[21][23] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2123_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3674_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2123_ ),
    .Y(\soc/cpu/cpuregs/_2124_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3675_  (.A0(\soc/cpu/cpuregs/regs[18][23] ),
    .A1(\soc/cpu/cpuregs/regs[19][23] ),
    .A2(\soc/cpu/cpuregs/regs[22][23] ),
    .A3(\soc/cpu/cpuregs/regs[23][23] ),
    .S0(net345),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2125_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3676_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2125_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2126_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3677_  (.A0(\soc/cpu/cpuregs/regs[2][23] ),
    .A1(\soc/cpu/cpuregs/regs[3][23] ),
    .A2(\soc/cpu/cpuregs/regs[6][23] ),
    .A3(\soc/cpu/cpuregs/regs[7][23] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2127_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3678_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2127_ ),
    .Y(\soc/cpu/cpuregs/_2128_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3679_  (.A0(\soc/cpu/cpuregs/regs[0][23] ),
    .A1(\soc/cpu/cpuregs/regs[1][23] ),
    .A2(\soc/cpu/cpuregs/regs[4][23] ),
    .A3(\soc/cpu/cpuregs/regs[5][23] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2129_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3680_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2129_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2130_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3681_  (.A1(\soc/cpu/cpuregs/_2124_ ),
    .A2(\soc/cpu/cpuregs/_2126_ ),
    .B1(\soc/cpu/cpuregs/_2128_ ),
    .B2(\soc/cpu/cpuregs/_2130_ ),
    .Y(\soc/cpu/cpuregs/_2131_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3682_  (.A0(\soc/cpu/cpuregs/regs[24][23] ),
    .A1(\soc/cpu/cpuregs/regs[25][23] ),
    .A2(\soc/cpu/cpuregs/regs[28][23] ),
    .A3(\soc/cpu/cpuregs/regs[29][23] ),
    .S0(net345),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2132_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3683_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2132_ ),
    .Y(\soc/cpu/cpuregs/_2133_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3684_  (.A0(\soc/cpu/cpuregs/regs[26][23] ),
    .A1(\soc/cpu/cpuregs/regs[27][23] ),
    .A2(\soc/cpu/cpuregs/regs[30][23] ),
    .A3(\soc/cpu/cpuregs/regs[31][23] ),
    .S0(net345),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2134_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3685_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2134_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2135_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3686_  (.A0(\soc/cpu/cpuregs/regs[10][23] ),
    .A1(\soc/cpu/cpuregs/regs[11][23] ),
    .A2(\soc/cpu/cpuregs/regs[14][23] ),
    .A3(\soc/cpu/cpuregs/regs[15][23] ),
    .S0(net345),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2136_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3687_  (.A0(\soc/cpu/cpuregs/regs[8][23] ),
    .A1(\soc/cpu/cpuregs/regs[9][23] ),
    .A2(\soc/cpu/cpuregs/regs[12][23] ),
    .A3(\soc/cpu/cpuregs/regs[13][23] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2137_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_3688_  (.A0(\soc/cpu/cpuregs/_2136_ ),
    .A1(\soc/cpu/cpuregs/_2137_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_2138_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3689_  (.A1(\soc/cpu/cpuregs/_2133_ ),
    .A2(\soc/cpu/cpuregs/_2135_ ),
    .B1(\soc/cpu/cpuregs/_2138_ ),
    .B2(net328),
    .C1(net330),
    .Y(\soc/cpu/cpuregs/_2139_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3690_  (.A1(net332),
    .A2(\soc/cpu/cpuregs/_2131_ ),
    .B1(\soc/cpu/cpuregs/_2139_ ),
    .X(\soc/cpu/cpuregs_rdata1[23] ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/cpuregs/_3691_  (.A(\soc/cpu/cpuregs/regs[18][24] ),
    .SLEEP(net338),
    .X(\soc/cpu/cpuregs/_2140_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/cpuregs/_3692_  (.A1(\soc/cpu/cpuregs/regs[22][24] ),
    .A2(net338),
    .B1(\soc/cpu/cpuregs/_2140_ ),
    .C1(net353),
    .X(\soc/cpu/cpuregs/_2141_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3693_  (.A0(\soc/cpu/cpuregs/regs[19][24] ),
    .A1(\soc/cpu/cpuregs/regs[23][24] ),
    .S(net338),
    .Y(\soc/cpu/cpuregs/_2142_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3694_  (.A1(net353),
    .A2(\soc/cpu/cpuregs/_2142_ ),
    .B1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_2143_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3695_  (.A0(\soc/cpu/cpuregs/regs[26][24] ),
    .A1(\soc/cpu/cpuregs/regs[27][24] ),
    .A2(\soc/cpu/cpuregs/regs[30][24] ),
    .A3(\soc/cpu/cpuregs/regs[31][24] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2144_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/cpuregs/_3696_  (.A1(\soc/cpu/cpuregs/_2141_ ),
    .A2(\soc/cpu/cpuregs/_2143_ ),
    .B1(\soc/cpu/cpuregs/_2144_ ),
    .B2(\soc/cpu/cpuregs_raddr1[3] ),
    .X(\soc/cpu/cpuregs/_2145_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3697_  (.A0(\soc/cpu/cpuregs/regs[16][24] ),
    .A1(\soc/cpu/cpuregs/regs[17][24] ),
    .A2(\soc/cpu/cpuregs/regs[20][24] ),
    .A3(\soc/cpu/cpuregs/regs[21][24] ),
    .S0(net353),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2146_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3698_  (.A0(\soc/cpu/cpuregs/regs[24][24] ),
    .A1(\soc/cpu/cpuregs/regs[25][24] ),
    .A2(\soc/cpu/cpuregs/regs[28][24] ),
    .A3(\soc/cpu/cpuregs/regs[29][24] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2147_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3699_  (.A0(\soc/cpu/cpuregs/_2146_ ),
    .A1(\soc/cpu/cpuregs/_2147_ ),
    .S(\soc/cpu/cpuregs_raddr1[3] ),
    .X(\soc/cpu/cpuregs/_2148_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3700_  (.A0(\soc/cpu/cpuregs/regs[10][24] ),
    .A1(\soc/cpu/cpuregs/regs[11][24] ),
    .A2(\soc/cpu/cpuregs/regs[14][24] ),
    .A3(\soc/cpu/cpuregs/regs[15][24] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2149_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/cpu/cpuregs/_3701_  (.A(\soc/cpu/cpuregs/regs[2][24] ),
    .SLEEP(net339),
    .X(\soc/cpu/cpuregs/_2150_ ));
 sky130_fd_sc_hd__a211o_1 \soc/cpu/cpuregs/_3702_  (.A1(\soc/cpu/cpuregs/regs[6][24] ),
    .A2(net339),
    .B1(\soc/cpu/cpuregs/_2150_ ),
    .C1(net353),
    .X(\soc/cpu/cpuregs/_2151_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3703_  (.A0(\soc/cpu/cpuregs/regs[3][24] ),
    .A1(\soc/cpu/cpuregs/regs[7][24] ),
    .S(net339),
    .Y(\soc/cpu/cpuregs/_2152_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3704_  (.A1(net353),
    .A2(\soc/cpu/cpuregs/_2152_ ),
    .B1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_2153_ ));
 sky130_fd_sc_hd__a22o_1 \soc/cpu/cpuregs/_3705_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_2149_ ),
    .B1(\soc/cpu/cpuregs/_2151_ ),
    .B2(\soc/cpu/cpuregs/_2153_ ),
    .X(\soc/cpu/cpuregs/_2154_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3706_  (.A0(\soc/cpu/cpuregs/regs[0][24] ),
    .A1(\soc/cpu/cpuregs/regs[1][24] ),
    .A2(\soc/cpu/cpuregs/regs[4][24] ),
    .A3(\soc/cpu/cpuregs/regs[5][24] ),
    .S0(net353),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2155_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3707_  (.A0(\soc/cpu/cpuregs/regs[8][24] ),
    .A1(\soc/cpu/cpuregs/regs[9][24] ),
    .A2(\soc/cpu/cpuregs/regs[12][24] ),
    .A3(\soc/cpu/cpuregs/regs[13][24] ),
    .S0(net352),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2156_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3708_  (.A0(\soc/cpu/cpuregs/_2155_ ),
    .A1(\soc/cpu/cpuregs/_2156_ ),
    .S(net332),
    .X(\soc/cpu/cpuregs/_2157_ ));
 sky130_fd_sc_hd__mux4_4 \soc/cpu/cpuregs/_3709_  (.A0(\soc/cpu/cpuregs/_2145_ ),
    .A1(\soc/cpu/cpuregs/_2148_ ),
    .A2(\soc/cpu/cpuregs/_2154_ ),
    .A3(\soc/cpu/cpuregs/_2157_ ),
    .S0(\soc/cpu/cpuregs/_1677_ ),
    .S1(\soc/cpu/cpuregs/_1699_ ),
    .X(\soc/cpu/cpuregs_rdata1[24] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3710_  (.A0(\soc/cpu/cpuregs/regs[16][25] ),
    .A1(\soc/cpu/cpuregs/regs[17][25] ),
    .A2(\soc/cpu/cpuregs/regs[20][25] ),
    .A3(\soc/cpu/cpuregs/regs[21][25] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2158_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3711_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2158_ ),
    .Y(\soc/cpu/cpuregs/_2159_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3712_  (.A0(\soc/cpu/cpuregs/regs[18][25] ),
    .A1(\soc/cpu/cpuregs/regs[19][25] ),
    .A2(\soc/cpu/cpuregs/regs[22][25] ),
    .A3(\soc/cpu/cpuregs/regs[23][25] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2160_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3713_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_2160_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_2161_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3714_  (.A0(\soc/cpu/cpuregs/regs[2][25] ),
    .A1(\soc/cpu/cpuregs/regs[3][25] ),
    .A2(\soc/cpu/cpuregs/regs[6][25] ),
    .A3(\soc/cpu/cpuregs/regs[7][25] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2162_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3715_  (.A(net152),
    .B(\soc/cpu/cpuregs/_2162_ ),
    .Y(\soc/cpu/cpuregs/_2163_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3716_  (.A0(\soc/cpu/cpuregs/regs[0][25] ),
    .A1(\soc/cpu/cpuregs/regs[1][25] ),
    .A2(\soc/cpu/cpuregs/regs[4][25] ),
    .A3(\soc/cpu/cpuregs/regs[5][25] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2164_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3717_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2164_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2165_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3718_  (.A1(\soc/cpu/cpuregs/_2159_ ),
    .A2(\soc/cpu/cpuregs/_2161_ ),
    .B1(\soc/cpu/cpuregs/_2163_ ),
    .B2(\soc/cpu/cpuregs/_2165_ ),
    .Y(\soc/cpu/cpuregs/_2166_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3719_  (.A0(\soc/cpu/cpuregs/regs[24][25] ),
    .A1(\soc/cpu/cpuregs/regs[25][25] ),
    .A2(\soc/cpu/cpuregs/regs[28][25] ),
    .A3(\soc/cpu/cpuregs/regs[29][25] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2167_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3720_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2167_ ),
    .Y(\soc/cpu/cpuregs/_2168_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3721_  (.A0(\soc/cpu/cpuregs/regs[26][25] ),
    .A1(\soc/cpu/cpuregs/regs[27][25] ),
    .A2(\soc/cpu/cpuregs/regs[30][25] ),
    .A3(\soc/cpu/cpuregs/regs[31][25] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2169_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3722_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_2169_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_2170_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3723_  (.A0(\soc/cpu/cpuregs/regs[10][25] ),
    .A1(\soc/cpu/cpuregs/regs[11][25] ),
    .A2(\soc/cpu/cpuregs/regs[14][25] ),
    .A3(\soc/cpu/cpuregs/regs[15][25] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2171_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3724_  (.A(net152),
    .B(\soc/cpu/cpuregs/_2171_ ),
    .Y(\soc/cpu/cpuregs/_2172_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3725_  (.A0(\soc/cpu/cpuregs/regs[8][25] ),
    .A1(\soc/cpu/cpuregs/regs[9][25] ),
    .A2(\soc/cpu/cpuregs/regs[12][25] ),
    .A3(\soc/cpu/cpuregs/regs[13][25] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2173_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3726_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2173_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2174_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3727_  (.A1(\soc/cpu/cpuregs/_2168_ ),
    .A2(\soc/cpu/cpuregs/_2170_ ),
    .B1(\soc/cpu/cpuregs/_2172_ ),
    .B2(\soc/cpu/cpuregs/_2174_ ),
    .C1(net332),
    .Y(\soc/cpu/cpuregs/_2175_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3728_  (.A1(net332),
    .A2(\soc/cpu/cpuregs/_2166_ ),
    .B1(\soc/cpu/cpuregs/_2175_ ),
    .X(\soc/cpu/cpuregs_rdata1[25] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3729_  (.A0(\soc/cpu/cpuregs/regs[16][26] ),
    .A1(\soc/cpu/cpuregs/regs[17][26] ),
    .A2(\soc/cpu/cpuregs/regs[20][26] ),
    .A3(\soc/cpu/cpuregs/regs[21][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2176_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3730_  (.A(net341),
    .B(\soc/cpu/cpuregs/_2176_ ),
    .Y(\soc/cpu/cpuregs/_2177_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3731_  (.A0(\soc/cpu/cpuregs/regs[18][26] ),
    .A1(\soc/cpu/cpuregs/regs[19][26] ),
    .A2(\soc/cpu/cpuregs/regs[22][26] ),
    .A3(\soc/cpu/cpuregs/regs[23][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2178_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3732_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2178_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2179_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3733_  (.A0(\soc/cpu/cpuregs/regs[2][26] ),
    .A1(\soc/cpu/cpuregs/regs[3][26] ),
    .A2(\soc/cpu/cpuregs/regs[6][26] ),
    .A3(\soc/cpu/cpuregs/regs[7][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2180_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3734_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2180_ ),
    .Y(\soc/cpu/cpuregs/_2181_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3735_  (.A0(\soc/cpu/cpuregs/regs[0][26] ),
    .A1(\soc/cpu/cpuregs/regs[1][26] ),
    .A2(\soc/cpu/cpuregs/regs[4][26] ),
    .A3(\soc/cpu/cpuregs/regs[5][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2182_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3736_  (.A1(net341),
    .A2(\soc/cpu/cpuregs/_2182_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2183_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3737_  (.A1(\soc/cpu/cpuregs/_2177_ ),
    .A2(\soc/cpu/cpuregs/_2179_ ),
    .B1(\soc/cpu/cpuregs/_2181_ ),
    .B2(\soc/cpu/cpuregs/_2183_ ),
    .Y(\soc/cpu/cpuregs/_2184_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3738_  (.A0(\soc/cpu/cpuregs/regs[24][26] ),
    .A1(\soc/cpu/cpuregs/regs[25][26] ),
    .A2(\soc/cpu/cpuregs/regs[28][26] ),
    .A3(\soc/cpu/cpuregs/regs[29][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2185_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3739_  (.A(net341),
    .B(\soc/cpu/cpuregs/_2185_ ),
    .Y(\soc/cpu/cpuregs/_2186_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3740_  (.A0(\soc/cpu/cpuregs/regs[26][26] ),
    .A1(\soc/cpu/cpuregs/regs[27][26] ),
    .A2(\soc/cpu/cpuregs/regs[30][26] ),
    .A3(\soc/cpu/cpuregs/regs[31][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2187_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3741_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2187_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2188_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3742_  (.A0(\soc/cpu/cpuregs/regs[10][26] ),
    .A1(\soc/cpu/cpuregs/regs[11][26] ),
    .A2(\soc/cpu/cpuregs/regs[14][26] ),
    .A3(\soc/cpu/cpuregs/regs[15][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2189_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3743_  (.A0(\soc/cpu/cpuregs/regs[8][26] ),
    .A1(\soc/cpu/cpuregs/regs[9][26] ),
    .A2(\soc/cpu/cpuregs/regs[12][26] ),
    .A3(\soc/cpu/cpuregs/regs[13][26] ),
    .S0(net347),
    .S1(net335),
    .X(\soc/cpu/cpuregs/_2190_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3744_  (.A0(\soc/cpu/cpuregs/_2189_ ),
    .A1(\soc/cpu/cpuregs/_2190_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2191_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3745_  (.A1(\soc/cpu/cpuregs/_2186_ ),
    .A2(\soc/cpu/cpuregs/_2188_ ),
    .B1(\soc/cpu/cpuregs/_2191_ ),
    .B2(net328),
    .C1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_2192_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/cpuregs/_3746_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_2184_ ),
    .B1(\soc/cpu/cpuregs/_2192_ ),
    .X(\soc/cpu/cpuregs_rdata1[26] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3747_  (.A0(\soc/cpu/cpuregs/regs[2][27] ),
    .A1(\soc/cpu/cpuregs/regs[3][27] ),
    .A2(\soc/cpu/cpuregs/regs[6][27] ),
    .A3(\soc/cpu/cpuregs/regs[7][27] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2193_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3748_  (.A0(\soc/cpu/cpuregs/regs[0][27] ),
    .A1(\soc/cpu/cpuregs/regs[1][27] ),
    .A2(\soc/cpu/cpuregs/regs[4][27] ),
    .A3(\soc/cpu/cpuregs/regs[5][27] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2194_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3749_  (.A0(\soc/cpu/cpuregs/_2193_ ),
    .A1(\soc/cpu/cpuregs/_2194_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_2195_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3750_  (.A0(\soc/cpu/cpuregs/regs[16][27] ),
    .A1(\soc/cpu/cpuregs/regs[17][27] ),
    .A2(\soc/cpu/cpuregs/regs[20][27] ),
    .A3(\soc/cpu/cpuregs/regs[21][27] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2196_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3751_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_2196_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2197_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3752_  (.A0(\soc/cpu/cpuregs/regs[18][27] ),
    .A1(\soc/cpu/cpuregs/regs[19][27] ),
    .A2(\soc/cpu/cpuregs/regs[22][27] ),
    .A3(\soc/cpu/cpuregs/regs[23][27] ),
    .S0(net345),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2198_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_3753_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2198_ ),
    .Y(\soc/cpu/cpuregs/_2199_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/cpuregs/_3754_  (.A1(\soc/cpu/cpuregs/_1699_ ),
    .A2(\soc/cpu/cpuregs/_2195_ ),
    .B1(\soc/cpu/cpuregs/_2197_ ),
    .B2(\soc/cpu/cpuregs/_2199_ ),
    .Y(\soc/cpu/cpuregs/_2200_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3755_  (.A0(\soc/cpu/cpuregs/regs[10][27] ),
    .A1(\soc/cpu/cpuregs/regs[11][27] ),
    .A2(\soc/cpu/cpuregs/regs[14][27] ),
    .A3(\soc/cpu/cpuregs/regs[15][27] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2201_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3756_  (.A0(\soc/cpu/cpuregs/regs[8][27] ),
    .A1(\soc/cpu/cpuregs/regs[9][27] ),
    .A2(\soc/cpu/cpuregs/regs[12][27] ),
    .A3(\soc/cpu/cpuregs/regs[13][27] ),
    .S0(net352),
    .S1(net337),
    .X(\soc/cpu/cpuregs/_2202_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_3757_  (.A0(\soc/cpu/cpuregs/_2201_ ),
    .A1(\soc/cpu/cpuregs/_2202_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_2203_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3758_  (.A0(\soc/cpu/cpuregs/regs[26][27] ),
    .A1(\soc/cpu/cpuregs/regs[27][27] ),
    .A2(\soc/cpu/cpuregs/regs[30][27] ),
    .A3(\soc/cpu/cpuregs/regs[31][27] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2204_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3759_  (.A(net152),
    .B(\soc/cpu/cpuregs/_2204_ ),
    .Y(\soc/cpu/cpuregs/_2205_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3760_  (.A0(\soc/cpu/cpuregs/regs[24][27] ),
    .A1(\soc/cpu/cpuregs/regs[25][27] ),
    .A2(\soc/cpu/cpuregs/regs[28][27] ),
    .A3(\soc/cpu/cpuregs/regs[29][27] ),
    .S0(net344),
    .S1(net333),
    .X(\soc/cpu/cpuregs/_2206_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3761_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2206_ ),
    .B1(net327),
    .Y(\soc/cpu/cpuregs/_2207_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3762_  (.A1(net327),
    .A2(\soc/cpu/cpuregs/_2203_ ),
    .B1(\soc/cpu/cpuregs/_2205_ ),
    .B2(\soc/cpu/cpuregs/_2207_ ),
    .C1(net332),
    .Y(\soc/cpu/cpuregs/_2208_ ));
 sky130_fd_sc_hd__o21a_2 \soc/cpu/cpuregs/_3763_  (.A1(net332),
    .A2(\soc/cpu/cpuregs/_2200_ ),
    .B1(\soc/cpu/cpuregs/_2208_ ),
    .X(\soc/cpu/cpuregs_rdata1[27] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3764_  (.A0(\soc/cpu/cpuregs/regs[16][28] ),
    .A1(\soc/cpu/cpuregs/regs[17][28] ),
    .A2(\soc/cpu/cpuregs/regs[20][28] ),
    .A3(\soc/cpu/cpuregs/regs[21][28] ),
    .S0(net348),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2209_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3765_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2209_ ),
    .Y(\soc/cpu/cpuregs/_2210_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3766_  (.A0(\soc/cpu/cpuregs/regs[18][28] ),
    .A1(\soc/cpu/cpuregs/regs[19][28] ),
    .A2(\soc/cpu/cpuregs/regs[22][28] ),
    .A3(\soc/cpu/cpuregs/regs[23][28] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2211_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3767_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2211_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2212_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3768_  (.A0(\soc/cpu/cpuregs/regs[2][28] ),
    .A1(\soc/cpu/cpuregs/regs[3][28] ),
    .A2(\soc/cpu/cpuregs/regs[6][28] ),
    .A3(\soc/cpu/cpuregs/regs[7][28] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2213_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3769_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2213_ ),
    .Y(\soc/cpu/cpuregs/_2214_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3770_  (.A0(\soc/cpu/cpuregs/regs[0][28] ),
    .A1(\soc/cpu/cpuregs/regs[1][28] ),
    .A2(\soc/cpu/cpuregs/regs[4][28] ),
    .A3(\soc/cpu/cpuregs/regs[5][28] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2215_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3771_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2215_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2216_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3772_  (.A1(\soc/cpu/cpuregs/_2210_ ),
    .A2(\soc/cpu/cpuregs/_2212_ ),
    .B1(\soc/cpu/cpuregs/_2214_ ),
    .B2(\soc/cpu/cpuregs/_2216_ ),
    .Y(\soc/cpu/cpuregs/_2217_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3773_  (.A0(\soc/cpu/cpuregs/regs[24][28] ),
    .A1(\soc/cpu/cpuregs/regs[25][28] ),
    .A2(\soc/cpu/cpuregs/regs[28][28] ),
    .A3(\soc/cpu/cpuregs/regs[29][28] ),
    .S0(net348),
    .S1(net334),
    .X(\soc/cpu/cpuregs/_2218_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3774_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2218_ ),
    .Y(\soc/cpu/cpuregs/_2219_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3775_  (.A0(\soc/cpu/cpuregs/regs[26][28] ),
    .A1(\soc/cpu/cpuregs/regs[27][28] ),
    .A2(\soc/cpu/cpuregs/regs[30][28] ),
    .A3(\soc/cpu/cpuregs/regs[31][28] ),
    .S0(net348),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2220_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3776_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2220_ ),
    .B1(net328),
    .Y(\soc/cpu/cpuregs/_2221_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3777_  (.A0(\soc/cpu/cpuregs/regs[10][28] ),
    .A1(\soc/cpu/cpuregs/regs[11][28] ),
    .A2(\soc/cpu/cpuregs/regs[14][28] ),
    .A3(\soc/cpu/cpuregs/regs[15][28] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2222_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3778_  (.A0(\soc/cpu/cpuregs/regs[8][28] ),
    .A1(\soc/cpu/cpuregs/regs[9][28] ),
    .A2(\soc/cpu/cpuregs/regs[12][28] ),
    .A3(\soc/cpu/cpuregs/regs[13][28] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2223_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3779_  (.A0(\soc/cpu/cpuregs/_2222_ ),
    .A1(\soc/cpu/cpuregs/_2223_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2224_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3780_  (.A1(\soc/cpu/cpuregs/_2219_ ),
    .A2(\soc/cpu/cpuregs/_2221_ ),
    .B1(\soc/cpu/cpuregs/_2224_ ),
    .B2(net328),
    .C1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_2225_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/cpuregs/_3781_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_2217_ ),
    .B1(\soc/cpu/cpuregs/_2225_ ),
    .X(\soc/cpu/cpuregs_rdata1[28] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3782_  (.A0(\soc/cpu/cpuregs/regs[16][29] ),
    .A1(\soc/cpu/cpuregs/regs[17][29] ),
    .A2(\soc/cpu/cpuregs/regs[20][29] ),
    .A3(\soc/cpu/cpuregs/regs[21][29] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2226_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3783_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2226_ ),
    .Y(\soc/cpu/cpuregs/_2227_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3784_  (.A0(\soc/cpu/cpuregs/regs[18][29] ),
    .A1(\soc/cpu/cpuregs/regs[19][29] ),
    .A2(\soc/cpu/cpuregs/regs[22][29] ),
    .A3(\soc/cpu/cpuregs/regs[23][29] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2228_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3785_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2228_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2229_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3786_  (.A0(\soc/cpu/cpuregs/regs[2][29] ),
    .A1(\soc/cpu/cpuregs/regs[3][29] ),
    .A2(\soc/cpu/cpuregs/regs[6][29] ),
    .A3(\soc/cpu/cpuregs/regs[7][29] ),
    .S0(net353),
    .S1(net340),
    .X(\soc/cpu/cpuregs/_2230_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3787_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2230_ ),
    .Y(\soc/cpu/cpuregs/_2231_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3788_  (.A0(\soc/cpu/cpuregs/regs[0][29] ),
    .A1(\soc/cpu/cpuregs/regs[1][29] ),
    .A2(\soc/cpu/cpuregs/regs[4][29] ),
    .A3(\soc/cpu/cpuregs/regs[5][29] ),
    .S0(net353),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2232_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3789_  (.A1(net343),
    .A2(\soc/cpu/cpuregs/_2232_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2233_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/cpu/cpuregs/_3790_  (.A1(\soc/cpu/cpuregs/_2227_ ),
    .A2(\soc/cpu/cpuregs/_2229_ ),
    .B1(\soc/cpu/cpuregs/_2231_ ),
    .B2(\soc/cpu/cpuregs/_2233_ ),
    .Y(\soc/cpu/cpuregs/_2234_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3791_  (.A0(\soc/cpu/cpuregs/regs[24][29] ),
    .A1(\soc/cpu/cpuregs/regs[25][29] ),
    .A2(\soc/cpu/cpuregs/regs[28][29] ),
    .A3(\soc/cpu/cpuregs/regs[29][29] ),
    .S0(net348),
    .S1(net336),
    .X(\soc/cpu/cpuregs/_2235_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3792_  (.A(net343),
    .B(\soc/cpu/cpuregs/_2235_ ),
    .Y(\soc/cpu/cpuregs/_2236_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3793_  (.A0(\soc/cpu/cpuregs/regs[26][29] ),
    .A1(\soc/cpu/cpuregs/regs[27][29] ),
    .A2(\soc/cpu/cpuregs/regs[30][29] ),
    .A3(\soc/cpu/cpuregs/regs[31][29] ),
    .S0(net348),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2237_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3794_  (.A1(\soc/cpu/cpuregs/_1677_ ),
    .A2(\soc/cpu/cpuregs/_2237_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2238_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3795_  (.A0(\soc/cpu/cpuregs/regs[10][29] ),
    .A1(\soc/cpu/cpuregs/regs[11][29] ),
    .A2(\soc/cpu/cpuregs/regs[14][29] ),
    .A3(\soc/cpu/cpuregs/regs[15][29] ),
    .S0(net353),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2239_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3796_  (.A0(\soc/cpu/cpuregs/regs[8][29] ),
    .A1(\soc/cpu/cpuregs/regs[9][29] ),
    .A2(\soc/cpu/cpuregs/regs[12][29] ),
    .A3(\soc/cpu/cpuregs/regs[13][29] ),
    .S0(net353),
    .S1(\soc/cpu/cpuregs_raddr1[2] ),
    .X(\soc/cpu/cpuregs/_2240_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3797_  (.A0(\soc/cpu/cpuregs/_2239_ ),
    .A1(\soc/cpu/cpuregs/_2240_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2241_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/cpu/cpuregs/_3798_  (.A1(\soc/cpu/cpuregs/_2236_ ),
    .A2(\soc/cpu/cpuregs/_2238_ ),
    .B1(\soc/cpu/cpuregs/_2241_ ),
    .B2(net329),
    .C1(\soc/cpu/cpuregs_raddr1[3] ),
    .Y(\soc/cpu/cpuregs/_2242_ ));
 sky130_fd_sc_hd__o21a_1 \soc/cpu/cpuregs/_3799_  (.A1(\soc/cpu/cpuregs_raddr1[3] ),
    .A2(\soc/cpu/cpuregs/_2234_ ),
    .B1(\soc/cpu/cpuregs/_2242_ ),
    .X(\soc/cpu/cpuregs_rdata1[29] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3800_  (.A0(\soc/cpu/cpuregs/regs[16][30] ),
    .A1(\soc/cpu/cpuregs/regs[17][30] ),
    .A2(\soc/cpu/cpuregs/regs[20][30] ),
    .A3(\soc/cpu/cpuregs/regs[21][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2243_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3801_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2243_ ),
    .Y(\soc/cpu/cpuregs/_2244_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3802_  (.A0(\soc/cpu/cpuregs/regs[18][30] ),
    .A1(\soc/cpu/cpuregs/regs[19][30] ),
    .A2(\soc/cpu/cpuregs/regs[22][30] ),
    .A3(\soc/cpu/cpuregs/regs[23][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2245_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3803_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_2245_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2246_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3804_  (.A0(\soc/cpu/cpuregs/regs[2][30] ),
    .A1(\soc/cpu/cpuregs/regs[3][30] ),
    .A2(\soc/cpu/cpuregs/regs[6][30] ),
    .A3(\soc/cpu/cpuregs/regs[7][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2247_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3805_  (.A(\soc/cpu/cpuregs/_1677_ ),
    .B(\soc/cpu/cpuregs/_2247_ ),
    .Y(\soc/cpu/cpuregs/_2248_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3806_  (.A0(\soc/cpu/cpuregs/regs[0][30] ),
    .A1(\soc/cpu/cpuregs/regs[1][30] ),
    .A2(\soc/cpu/cpuregs/regs[4][30] ),
    .A3(\soc/cpu/cpuregs/regs[5][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2249_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/cpu/cpuregs/_3807_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_2249_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2250_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/cpu/cpuregs/_3808_  (.A1(\soc/cpu/cpuregs/_2244_ ),
    .A2(\soc/cpu/cpuregs/_2246_ ),
    .B1(\soc/cpu/cpuregs/_2248_ ),
    .B2(\soc/cpu/cpuregs/_2250_ ),
    .Y(\soc/cpu/cpuregs/_2251_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3809_  (.A0(\soc/cpu/cpuregs/regs[24][30] ),
    .A1(\soc/cpu/cpuregs/regs[25][30] ),
    .A2(\soc/cpu/cpuregs/regs[28][30] ),
    .A3(\soc/cpu/cpuregs/regs[29][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2252_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3810_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2252_ ),
    .Y(\soc/cpu/cpuregs/_2253_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3811_  (.A0(\soc/cpu/cpuregs/regs[26][30] ),
    .A1(\soc/cpu/cpuregs/regs[27][30] ),
    .A2(\soc/cpu/cpuregs/regs[30][30] ),
    .A3(\soc/cpu/cpuregs/regs[31][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2254_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3812_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_2254_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2255_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3813_  (.A0(\soc/cpu/cpuregs/regs[10][30] ),
    .A1(\soc/cpu/cpuregs/regs[11][30] ),
    .A2(\soc/cpu/cpuregs/regs[14][30] ),
    .A3(\soc/cpu/cpuregs/regs[15][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2256_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3814_  (.A0(\soc/cpu/cpuregs/regs[8][30] ),
    .A1(\soc/cpu/cpuregs/regs[9][30] ),
    .A2(\soc/cpu/cpuregs/regs[12][30] ),
    .A3(\soc/cpu/cpuregs/regs[13][30] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2257_ ));
 sky130_fd_sc_hd__mux2i_2 \soc/cpu/cpuregs/_3815_  (.A0(\soc/cpu/cpuregs/_2256_ ),
    .A1(\soc/cpu/cpuregs/_2257_ ),
    .S(\soc/cpu/cpuregs/_1677_ ),
    .Y(\soc/cpu/cpuregs/_2258_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/cpu/cpuregs/_3816_  (.A1(\soc/cpu/cpuregs/_2253_ ),
    .A2(\soc/cpu/cpuregs/_2255_ ),
    .B1(\soc/cpu/cpuregs/_2258_ ),
    .B2(net329),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_2259_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3817_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_2251_ ),
    .B1(\soc/cpu/cpuregs/_2259_ ),
    .X(\soc/cpu/cpuregs_rdata1[30] ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3818_  (.A0(\soc/cpu/cpuregs/regs[2][31] ),
    .A1(\soc/cpu/cpuregs/regs[3][31] ),
    .A2(\soc/cpu/cpuregs/regs[6][31] ),
    .A3(\soc/cpu/cpuregs/regs[7][31] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2260_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3819_  (.A0(\soc/cpu/cpuregs/regs[0][31] ),
    .A1(\soc/cpu/cpuregs/regs[1][31] ),
    .A2(\soc/cpu/cpuregs/regs[4][31] ),
    .A3(\soc/cpu/cpuregs/regs[5][31] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2261_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/cpu/cpuregs/_3820_  (.A0(\soc/cpu/cpuregs/_2260_ ),
    .A1(\soc/cpu/cpuregs/_2261_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_2262_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3821_  (.A0(\soc/cpu/cpuregs/regs[16][31] ),
    .A1(\soc/cpu/cpuregs/regs[17][31] ),
    .A2(\soc/cpu/cpuregs/regs[20][31] ),
    .A3(\soc/cpu/cpuregs/regs[21][31] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2263_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/cpu/cpuregs/_3822_  (.A1(net152),
    .A2(\soc/cpu/cpuregs/_2263_ ),
    .B1(\soc/cpu/cpuregs/_1699_ ),
    .Y(\soc/cpu/cpuregs/_2264_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3823_  (.A0(\soc/cpu/cpuregs/regs[18][31] ),
    .A1(\soc/cpu/cpuregs/regs[19][31] ),
    .A2(\soc/cpu/cpuregs/regs[22][31] ),
    .A3(\soc/cpu/cpuregs/regs[23][31] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2265_ ));
 sky130_fd_sc_hd__nand2_1 \soc/cpu/cpuregs/_3824_  (.A(net342),
    .B(\soc/cpu/cpuregs/_2265_ ),
    .Y(\soc/cpu/cpuregs/_2266_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/cpu/cpuregs/_3825_  (.A1(\soc/cpu/cpuregs/_1699_ ),
    .A2(\soc/cpu/cpuregs/_2262_ ),
    .B1(\soc/cpu/cpuregs/_2264_ ),
    .B2(\soc/cpu/cpuregs/_2266_ ),
    .Y(\soc/cpu/cpuregs/_2267_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3826_  (.A0(\soc/cpu/cpuregs/regs[10][31] ),
    .A1(\soc/cpu/cpuregs/regs[11][31] ),
    .A2(\soc/cpu/cpuregs/regs[14][31] ),
    .A3(\soc/cpu/cpuregs/regs[15][31] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2268_ ));
 sky130_fd_sc_hd__mux4_2 \soc/cpu/cpuregs/_3827_  (.A0(\soc/cpu/cpuregs/regs[8][31] ),
    .A1(\soc/cpu/cpuregs/regs[9][31] ),
    .A2(\soc/cpu/cpuregs/regs[12][31] ),
    .A3(\soc/cpu/cpuregs/regs[13][31] ),
    .S0(net349),
    .S1(net339),
    .X(\soc/cpu/cpuregs/_2269_ ));
 sky130_fd_sc_hd__mux2i_4 \soc/cpu/cpuregs/_3828_  (.A0(\soc/cpu/cpuregs/_2268_ ),
    .A1(\soc/cpu/cpuregs/_2269_ ),
    .S(net152),
    .Y(\soc/cpu/cpuregs/_2270_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3829_  (.A0(\soc/cpu/cpuregs/regs[26][31] ),
    .A1(\soc/cpu/cpuregs/regs[27][31] ),
    .A2(\soc/cpu/cpuregs/regs[30][31] ),
    .A3(\soc/cpu/cpuregs/regs[31][31] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2271_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_3830_  (.A(net152),
    .B(\soc/cpu/cpuregs/_2271_ ),
    .Y(\soc/cpu/cpuregs/_2272_ ));
 sky130_fd_sc_hd__mux4_1 \soc/cpu/cpuregs/_3831_  (.A0(\soc/cpu/cpuregs/regs[24][31] ),
    .A1(\soc/cpu/cpuregs/regs[25][31] ),
    .A2(\soc/cpu/cpuregs/regs[28][31] ),
    .A3(\soc/cpu/cpuregs/regs[29][31] ),
    .S0(net351),
    .S1(net338),
    .X(\soc/cpu/cpuregs/_2273_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/cpu/cpuregs/_3832_  (.A1(net342),
    .A2(\soc/cpu/cpuregs/_2273_ ),
    .B1(net329),
    .Y(\soc/cpu/cpuregs/_2274_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/cpu/cpuregs/_3833_  (.A1(net329),
    .A2(\soc/cpu/cpuregs/_2270_ ),
    .B1(\soc/cpu/cpuregs/_2272_ ),
    .B2(\soc/cpu/cpuregs/_2274_ ),
    .C1(net331),
    .Y(\soc/cpu/cpuregs/_2275_ ));
 sky130_fd_sc_hd__o21a_4 \soc/cpu/cpuregs/_3834_  (.A1(net331),
    .A2(\soc/cpu/cpuregs/_2267_ ),
    .B1(\soc/cpu/cpuregs/_2275_ ),
    .X(\soc/cpu/cpuregs_rdata1[31] ));
 sky130_fd_sc_hd__nand3b_4 \soc/cpu/cpuregs/_3836_  (.A_N(\soc/cpu/cpuregs_waddr[2] ),
    .B(\soc/cpu/cpuregs_waddr[3] ),
    .C(\soc/cpu/cpuregs_waddr[4] ),
    .Y(\soc/cpu/cpuregs/_2277_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/cpuregs/_3837_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/cpuregs_waddr[0] ),
    .C(\soc/cpu/_00074_ ),
    .Y(\soc/cpu/cpuregs/_2278_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_3838_  (.A(\soc/cpu/cpuregs/_2277_ ),
    .B(\soc/cpu/cpuregs/_2278_ ),
    .Y(\soc/cpu/cpuregs/_2279_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3840_  (.A0(\soc/cpu/cpuregs/regs[27][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0000_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3842_  (.A0(\soc/cpu/cpuregs/regs[27][1] ),
    .A1(net130),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0001_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3844_  (.A0(\soc/cpu/cpuregs/regs[27][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0002_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3846_  (.A0(\soc/cpu/cpuregs/regs[27][3] ),
    .A1(net129),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0003_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3848_  (.A0(\soc/cpu/cpuregs/regs[27][4] ),
    .A1(net128),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0004_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3850_  (.A0(\soc/cpu/cpuregs/regs[27][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0005_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3852_  (.A0(\soc/cpu/cpuregs/regs[27][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0006_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3854_  (.A0(\soc/cpu/cpuregs/regs[27][7] ),
    .A1(net125),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0007_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3856_  (.A0(\soc/cpu/cpuregs/regs[27][8] ),
    .A1(net127),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0008_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3858_  (.A0(\soc/cpu/cpuregs/regs[27][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0009_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3861_  (.A0(\soc/cpu/cpuregs/regs[27][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0010_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3863_  (.A0(\soc/cpu/cpuregs/regs[27][11] ),
    .A1(net124),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0011_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3865_  (.A0(\soc/cpu/cpuregs/regs[27][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0012_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3867_  (.A0(\soc/cpu/cpuregs/regs[27][13] ),
    .A1(net105),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0013_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3869_  (.A0(\soc/cpu/cpuregs/regs[27][14] ),
    .A1(net114),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0014_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3871_  (.A0(\soc/cpu/cpuregs/regs[27][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0015_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3873_  (.A0(\soc/cpu/cpuregs/regs[27][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0016_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3875_  (.A0(\soc/cpu/cpuregs/regs[27][17] ),
    .A1(net88),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0017_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3877_  (.A0(\soc/cpu/cpuregs/regs[27][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0018_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3879_  (.A0(\soc/cpu/cpuregs/regs[27][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0019_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3882_  (.A0(\soc/cpu/cpuregs/regs[27][20] ),
    .A1(net63),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0020_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3884_  (.A0(\soc/cpu/cpuregs/regs[27][21] ),
    .A1(net59),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0021_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3886_  (.A0(\soc/cpu/cpuregs/regs[27][22] ),
    .A1(net60),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0022_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3888_  (.A0(\soc/cpu/cpuregs/regs[27][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0023_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3890_  (.A0(\soc/cpu/cpuregs/regs[27][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0024_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3892_  (.A0(\soc/cpu/cpuregs/regs[27][25] ),
    .A1(net58),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0025_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3894_  (.A0(\soc/cpu/cpuregs/regs[27][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net103),
    .X(\soc/cpu/cpuregs/_0026_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3896_  (.A0(\soc/cpu/cpuregs/regs[27][27] ),
    .A1(net55),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0027_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3898_  (.A0(\soc/cpu/cpuregs/regs[27][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(\soc/cpu/cpuregs/_2279_ ),
    .X(\soc/cpu/cpuregs/_0028_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3900_  (.A0(\soc/cpu/cpuregs/regs[27][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0029_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3902_  (.A0(\soc/cpu/cpuregs/regs[27][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0030_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3904_  (.A0(\soc/cpu/cpuregs/regs[27][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net104),
    .X(\soc/cpu/cpuregs/_0031_ ));
 sky130_fd_sc_hd__nor3b_4 \soc/cpu/cpuregs/_3906_  (.A(\soc/cpu/cpuregs_waddr[3] ),
    .B(\soc/cpu/cpuregs_waddr[4] ),
    .C_N(\soc/cpu/cpuregs_waddr[2] ),
    .Y(\soc/cpu/cpuregs/_2315_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/cpuregs/_3907_  (.A(\soc/cpu/cpuregs_waddr[0] ),
    .B(\soc/cpu/_00074_ ),
    .Y(\soc/cpu/cpuregs/_2316_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_3908_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/cpuregs/_2316_ ),
    .Y(\soc/cpu/cpuregs/_2317_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_3909_  (.A(\soc/cpu/cpuregs/_2315_ ),
    .B(\soc/cpu/cpuregs/_2317_ ),
    .Y(\soc/cpu/cpuregs/_2318_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3911_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[5][0] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0032_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3913_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[5][1] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0033_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3915_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[5][2] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0034_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3917_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[5][3] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0035_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3919_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[5][4] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0036_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3921_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[5][5] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0037_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3923_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[5][6] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0038_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3925_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[5][7] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0039_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3927_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[5][8] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0040_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3929_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[5][9] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0041_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3932_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[5][10] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0042_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3934_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[5][11] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0043_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3936_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[5][12] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0044_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3938_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[5][13] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0045_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3940_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[5][14] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0046_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3942_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[5][15] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0047_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3944_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[5][16] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0048_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3946_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[5][17] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0049_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3948_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[5][18] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0050_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3950_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[5][19] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0051_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3953_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[5][20] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0052_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3955_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[5][21] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0053_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3957_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[5][22] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0054_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3959_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[5][23] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0055_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3961_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[5][24] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0056_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3963_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[5][25] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0057_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3965_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[5][26] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0058_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3967_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[5][27] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0059_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3969_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[5][28] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0060_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3971_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[5][29] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0061_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3973_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[5][30] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0062_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3975_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[5][31] ),
    .S(\soc/cpu/cpuregs/_2318_ ),
    .X(\soc/cpu/cpuregs/_0063_ ));
 sky130_fd_sc_hd__nand2_2 \soc/cpu/cpuregs/_3976_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/_00074_ ),
    .Y(\soc/cpu/cpuregs/_2353_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_3977_  (.A(\soc/cpu/cpuregs_waddr[0] ),
    .B(\soc/cpu/cpuregs/_2353_ ),
    .Y(\soc/cpu/cpuregs/_2354_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_3978_  (.A(\soc/cpu/cpuregs/_2315_ ),
    .B(\soc/cpu/cpuregs/_2354_ ),
    .Y(\soc/cpu/cpuregs/_2355_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3980_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[6][0] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0064_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3981_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[6][1] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0065_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3982_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[6][2] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0066_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3983_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[6][3] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0067_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3984_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[6][4] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0068_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3985_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[6][5] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0069_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3986_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[6][6] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0070_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3987_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[6][7] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0071_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3988_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[6][8] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0072_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3989_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[6][9] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0073_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3991_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[6][10] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0074_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3992_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[6][11] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0075_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3993_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[6][12] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0076_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3994_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[6][13] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0077_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3995_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[6][14] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0078_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3996_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[6][15] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0079_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3997_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[6][16] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0080_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3998_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[6][17] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0081_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_3999_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[6][18] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0082_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4000_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[6][19] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0083_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4002_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[6][20] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0084_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4003_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[6][21] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0085_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4004_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[6][22] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0086_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4005_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[6][23] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0087_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4006_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[6][24] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0088_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4007_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[6][25] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0089_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4008_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[6][26] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0090_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4009_  (.A0(net55),
    .A1(\soc/cpu/cpuregs/regs[6][27] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0091_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4010_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[6][28] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0092_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4011_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[6][29] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0093_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4012_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[6][30] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0094_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4013_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[6][31] ),
    .S(\soc/cpu/cpuregs/_2355_ ),
    .X(\soc/cpu/cpuregs/_0095_ ));
 sky130_fd_sc_hd__nand3b_4 \soc/cpu/cpuregs/_4014_  (.A_N(\soc/cpu/cpuregs_waddr[4] ),
    .B(\soc/cpu/cpuregs_waddr[3] ),
    .C(\soc/cpu/cpuregs_waddr[2] ),
    .Y(\soc/cpu/cpuregs/_2359_ ));
 sky130_fd_sc_hd__nor2_2 \soc/cpu/cpuregs/_4015_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/cpuregs_waddr[0] ),
    .Y(\soc/cpu/cpuregs/_2360_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4016_  (.A(\soc/cpu/_00074_ ),
    .B(\soc/cpu/cpuregs/_2360_ ),
    .Y(\soc/cpu/cpuregs/_2361_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4017_  (.A(\soc/cpu/cpuregs/_2359_ ),
    .B(\soc/cpu/cpuregs/_2361_ ),
    .Y(\soc/cpu/cpuregs/_2362_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4019_  (.A0(\soc/cpu/cpuregs/regs[12][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0096_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4020_  (.A0(\soc/cpu/cpuregs/regs[12][1] ),
    .A1(net130),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0097_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4021_  (.A0(\soc/cpu/cpuregs/regs[12][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0098_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4022_  (.A0(\soc/cpu/cpuregs/regs[12][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0099_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4023_  (.A0(\soc/cpu/cpuregs/regs[12][4] ),
    .A1(net128),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0100_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4024_  (.A0(\soc/cpu/cpuregs/regs[12][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0101_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4025_  (.A0(\soc/cpu/cpuregs/regs[12][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0102_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4026_  (.A0(\soc/cpu/cpuregs/regs[12][7] ),
    .A1(net125),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0103_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4027_  (.A0(\soc/cpu/cpuregs/regs[12][8] ),
    .A1(net126),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0104_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4028_  (.A0(\soc/cpu/cpuregs/regs[12][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0105_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4030_  (.A0(\soc/cpu/cpuregs/regs[12][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0106_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4031_  (.A0(\soc/cpu/cpuregs/regs[12][11] ),
    .A1(net124),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0107_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4032_  (.A0(\soc/cpu/cpuregs/regs[12][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0108_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4033_  (.A0(\soc/cpu/cpuregs/regs[12][13] ),
    .A1(net105),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0109_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4034_  (.A0(\soc/cpu/cpuregs/regs[12][14] ),
    .A1(net113),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0110_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4035_  (.A0(\soc/cpu/cpuregs/regs[12][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0111_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4036_  (.A0(\soc/cpu/cpuregs/regs[12][16] ),
    .A1(net69),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0112_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4037_  (.A0(\soc/cpu/cpuregs/regs[12][17] ),
    .A1(net87),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0113_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4038_  (.A0(\soc/cpu/cpuregs/regs[12][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0114_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4039_  (.A0(\soc/cpu/cpuregs/regs[12][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0115_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4041_  (.A0(\soc/cpu/cpuregs/regs[12][20] ),
    .A1(net63),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0116_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4042_  (.A0(\soc/cpu/cpuregs/regs[12][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0117_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4043_  (.A0(\soc/cpu/cpuregs/regs[12][22] ),
    .A1(net61),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0118_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4044_  (.A0(\soc/cpu/cpuregs/regs[12][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0119_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4045_  (.A0(\soc/cpu/cpuregs/regs[12][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0120_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4046_  (.A0(\soc/cpu/cpuregs/regs[12][25] ),
    .A1(net57),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0121_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4047_  (.A0(\soc/cpu/cpuregs/regs[12][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0122_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4048_  (.A0(\soc/cpu/cpuregs/regs[12][27] ),
    .A1(net56),
    .S(net102),
    .X(\soc/cpu/cpuregs/_0123_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4049_  (.A0(\soc/cpu/cpuregs/regs[12][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net101),
    .X(\soc/cpu/cpuregs/_0124_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4050_  (.A0(\soc/cpu/cpuregs/regs[12][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0125_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4051_  (.A0(\soc/cpu/cpuregs/regs[12][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0126_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4052_  (.A0(\soc/cpu/cpuregs/regs[12][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(\soc/cpu/cpuregs/_2362_ ),
    .X(\soc/cpu/cpuregs/_0127_ ));
 sky130_fd_sc_hd__nor3_4 \soc/cpu/cpuregs/_4053_  (.A(\soc/cpu/cpuregs_waddr[2] ),
    .B(\soc/cpu/cpuregs_waddr[3] ),
    .C(\soc/cpu/cpuregs_waddr[4] ),
    .Y(\soc/cpu/cpuregs/_2366_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4054_  (.A(\soc/cpu/cpuregs/_2317_ ),
    .B(\soc/cpu/cpuregs/_2366_ ),
    .Y(\soc/cpu/cpuregs/_2367_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4056_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[1][0] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0128_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4057_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[1][1] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0129_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4058_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[1][2] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0130_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4059_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[1][3] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0131_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4060_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[1][4] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0132_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4061_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[1][5] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0133_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4062_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[1][6] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0134_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4063_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[1][7] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0135_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4064_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[1][8] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0136_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4065_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[1][9] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0137_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4067_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[1][10] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0138_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4068_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[1][11] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0139_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4069_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[1][12] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0140_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4070_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[1][13] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0141_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4071_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[1][14] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0142_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4072_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[1][15] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0143_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4073_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[1][16] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0144_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4074_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[1][17] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0145_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4075_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[1][18] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0146_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4076_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[1][19] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0147_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4078_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[1][20] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0148_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4079_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[1][21] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0149_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4080_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[1][22] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0150_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4081_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[1][23] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0151_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4082_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[1][24] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0152_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4083_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[1][25] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0153_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4084_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[1][26] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0154_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4085_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[1][27] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0155_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4086_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[1][28] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0156_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4087_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[1][29] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0157_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4088_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[1][30] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0158_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4089_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[1][31] ),
    .S(\soc/cpu/cpuregs/_2367_ ),
    .X(\soc/cpu/cpuregs/_0159_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/cpuregs/_4090_  (.A(\soc/cpu/cpuregs_waddr[0] ),
    .B(\soc/cpu/cpuregs/_2353_ ),
    .X(\soc/cpu/cpuregs/_2371_ ));
 sky130_fd_sc_hd__nand3b_4 \soc/cpu/cpuregs/_4091_  (.A_N(\soc/cpu/cpuregs_waddr[3] ),
    .B(\soc/cpu/cpuregs_waddr[4] ),
    .C(\soc/cpu/cpuregs_waddr[2] ),
    .Y(\soc/cpu/cpuregs/_2372_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4092_  (.A(\soc/cpu/cpuregs/_2371_ ),
    .B(\soc/cpu/cpuregs/_2372_ ),
    .Y(\soc/cpu/cpuregs/_2373_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4094_  (.A0(\soc/cpu/cpuregs/regs[22][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0160_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4095_  (.A0(\soc/cpu/cpuregs/regs[22][1] ),
    .A1(net130),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0161_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4096_  (.A0(\soc/cpu/cpuregs/regs[22][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0162_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4097_  (.A0(\soc/cpu/cpuregs/regs[22][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0163_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4098_  (.A0(\soc/cpu/cpuregs/regs[22][4] ),
    .A1(net128),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0164_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4099_  (.A0(\soc/cpu/cpuregs/regs[22][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0165_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4100_  (.A0(\soc/cpu/cpuregs/regs[22][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0166_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4101_  (.A0(\soc/cpu/cpuregs/regs[22][7] ),
    .A1(net125),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0167_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4102_  (.A0(\soc/cpu/cpuregs/regs[22][8] ),
    .A1(net127),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0168_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4103_  (.A0(\soc/cpu/cpuregs/regs[22][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0169_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4105_  (.A0(\soc/cpu/cpuregs/regs[22][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0170_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4106_  (.A0(\soc/cpu/cpuregs/regs[22][11] ),
    .A1(net123),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0171_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4107_  (.A0(\soc/cpu/cpuregs/regs[22][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0172_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4108_  (.A0(\soc/cpu/cpuregs/regs[22][13] ),
    .A1(net105),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0173_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4109_  (.A0(\soc/cpu/cpuregs/regs[22][14] ),
    .A1(net113),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0174_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4110_  (.A0(\soc/cpu/cpuregs/regs[22][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0175_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4111_  (.A0(\soc/cpu/cpuregs/regs[22][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0176_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4112_  (.A0(\soc/cpu/cpuregs/regs[22][17] ),
    .A1(net88),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0177_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4113_  (.A0(\soc/cpu/cpuregs/regs[22][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0178_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4114_  (.A0(\soc/cpu/cpuregs/regs[22][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0179_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4116_  (.A0(\soc/cpu/cpuregs/regs[22][20] ),
    .A1(net64),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0180_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4117_  (.A0(\soc/cpu/cpuregs/regs[22][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0181_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4118_  (.A0(\soc/cpu/cpuregs/regs[22][22] ),
    .A1(net60),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0182_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4119_  (.A0(\soc/cpu/cpuregs/regs[22][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0183_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4120_  (.A0(\soc/cpu/cpuregs/regs[22][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0184_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4121_  (.A0(\soc/cpu/cpuregs/regs[22][25] ),
    .A1(net58),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0185_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4122_  (.A0(\soc/cpu/cpuregs/regs[22][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net85),
    .X(\soc/cpu/cpuregs/_0186_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4123_  (.A0(\soc/cpu/cpuregs/regs[22][27] ),
    .A1(net55),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0187_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4124_  (.A0(\soc/cpu/cpuregs/regs[22][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0188_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4125_  (.A0(\soc/cpu/cpuregs/regs[22][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0189_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4126_  (.A0(\soc/cpu/cpuregs/regs[22][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2373_ ),
    .X(\soc/cpu/cpuregs/_0190_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4127_  (.A0(\soc/cpu/cpuregs/regs[22][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net86),
    .X(\soc/cpu/cpuregs/_0191_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4128_  (.A(\soc/cpu/cpuregs/_2278_ ),
    .B(\soc/cpu/cpuregs/_2372_ ),
    .Y(\soc/cpu/cpuregs/_2377_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4130_  (.A0(\soc/cpu/cpuregs/regs[23][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0192_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4131_  (.A0(\soc/cpu/cpuregs/regs[23][1] ),
    .A1(net130),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0193_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4132_  (.A0(\soc/cpu/cpuregs/regs[23][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0194_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4133_  (.A0(\soc/cpu/cpuregs/regs[23][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0195_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4134_  (.A0(\soc/cpu/cpuregs/regs[23][4] ),
    .A1(net128),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0196_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4135_  (.A0(\soc/cpu/cpuregs/regs[23][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0197_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4136_  (.A0(\soc/cpu/cpuregs/regs[23][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0198_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4137_  (.A0(\soc/cpu/cpuregs/regs[23][7] ),
    .A1(net125),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0199_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4138_  (.A0(\soc/cpu/cpuregs/regs[23][8] ),
    .A1(net127),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0200_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4139_  (.A0(\soc/cpu/cpuregs/regs[23][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0201_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4141_  (.A0(\soc/cpu/cpuregs/regs[23][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0202_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4142_  (.A0(\soc/cpu/cpuregs/regs[23][11] ),
    .A1(net123),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0203_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4143_  (.A0(\soc/cpu/cpuregs/regs[23][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0204_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4144_  (.A0(\soc/cpu/cpuregs/regs[23][13] ),
    .A1(net105),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0205_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4145_  (.A0(\soc/cpu/cpuregs/regs[23][14] ),
    .A1(net113),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0206_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4146_  (.A0(\soc/cpu/cpuregs/regs[23][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0207_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4147_  (.A0(\soc/cpu/cpuregs/regs[23][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0208_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4148_  (.A0(\soc/cpu/cpuregs/regs[23][17] ),
    .A1(net88),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0209_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4149_  (.A0(\soc/cpu/cpuregs/regs[23][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0210_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4150_  (.A0(\soc/cpu/cpuregs/regs[23][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0211_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4152_  (.A0(\soc/cpu/cpuregs/regs[23][20] ),
    .A1(net64),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0212_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4153_  (.A0(\soc/cpu/cpuregs/regs[23][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0213_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4154_  (.A0(\soc/cpu/cpuregs/regs[23][22] ),
    .A1(net60),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0214_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4155_  (.A0(\soc/cpu/cpuregs/regs[23][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0215_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4156_  (.A0(\soc/cpu/cpuregs/regs[23][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0216_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4157_  (.A0(\soc/cpu/cpuregs/regs[23][25] ),
    .A1(net58),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0217_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4158_  (.A0(\soc/cpu/cpuregs/regs[23][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net99),
    .X(\soc/cpu/cpuregs/_0218_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4159_  (.A0(\soc/cpu/cpuregs/regs[23][27] ),
    .A1(net55),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0219_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4160_  (.A0(\soc/cpu/cpuregs/regs[23][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0220_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4161_  (.A0(\soc/cpu/cpuregs/regs[23][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0221_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4162_  (.A0(\soc/cpu/cpuregs/regs[23][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2377_ ),
    .X(\soc/cpu/cpuregs/_0222_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4163_  (.A0(\soc/cpu/cpuregs/regs[23][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net100),
    .X(\soc/cpu/cpuregs/_0223_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4165_  (.A(\soc/cpu/cpuregs/_2361_ ),
    .B(\soc/cpu/cpuregs/_2372_ ),
    .Y(\soc/cpu/cpuregs/_2382_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4167_  (.A0(\soc/cpu/cpuregs/regs[20][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0224_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4169_  (.A0(\soc/cpu/cpuregs/regs[20][1] ),
    .A1(net130),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0225_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4171_  (.A0(\soc/cpu/cpuregs/regs[20][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0226_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4173_  (.A0(\soc/cpu/cpuregs/regs[20][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0227_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4175_  (.A0(\soc/cpu/cpuregs/regs[20][4] ),
    .A1(net128),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0228_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4177_  (.A0(\soc/cpu/cpuregs/regs[20][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0229_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4179_  (.A0(\soc/cpu/cpuregs/regs[20][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0230_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4181_  (.A0(\soc/cpu/cpuregs/regs[20][7] ),
    .A1(net125),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0231_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4183_  (.A0(\soc/cpu/cpuregs/regs[20][8] ),
    .A1(net126),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0232_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4185_  (.A0(\soc/cpu/cpuregs/regs[20][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0233_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4188_  (.A0(\soc/cpu/cpuregs/regs[20][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0234_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4190_  (.A0(\soc/cpu/cpuregs/regs[20][11] ),
    .A1(net123),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0235_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4192_  (.A0(\soc/cpu/cpuregs/regs[20][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0236_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4194_  (.A0(\soc/cpu/cpuregs/regs[20][13] ),
    .A1(net105),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0237_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4196_  (.A0(\soc/cpu/cpuregs/regs[20][14] ),
    .A1(net113),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0238_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4198_  (.A0(\soc/cpu/cpuregs/regs[20][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0239_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4200_  (.A0(\soc/cpu/cpuregs/regs[20][16] ),
    .A1(net69),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0240_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4202_  (.A0(\soc/cpu/cpuregs/regs[20][17] ),
    .A1(net87),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0241_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4204_  (.A0(\soc/cpu/cpuregs/regs[20][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0242_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4206_  (.A0(\soc/cpu/cpuregs/regs[20][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0243_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4209_  (.A0(\soc/cpu/cpuregs/regs[20][20] ),
    .A1(net64),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0244_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4211_  (.A0(\soc/cpu/cpuregs/regs[20][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0245_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4213_  (.A0(\soc/cpu/cpuregs/regs[20][22] ),
    .A1(net61),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0246_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4215_  (.A0(\soc/cpu/cpuregs/regs[20][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0247_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4217_  (.A0(\soc/cpu/cpuregs/regs[20][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0248_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4219_  (.A0(\soc/cpu/cpuregs/regs[20][25] ),
    .A1(net57),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0249_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4221_  (.A0(\soc/cpu/cpuregs/regs[20][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0250_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4223_  (.A0(\soc/cpu/cpuregs/regs[20][27] ),
    .A1(net55),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0251_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4225_  (.A0(\soc/cpu/cpuregs/regs[20][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net98),
    .X(\soc/cpu/cpuregs/_0252_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4227_  (.A0(\soc/cpu/cpuregs/regs[20][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0253_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4229_  (.A0(\soc/cpu/cpuregs/regs[20][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2382_ ),
    .X(\soc/cpu/cpuregs/_0254_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4231_  (.A0(\soc/cpu/cpuregs/regs[20][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net97),
    .X(\soc/cpu/cpuregs/_0255_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4232_  (.A(\soc/cpu/cpuregs/_2277_ ),
    .B(\soc/cpu/cpuregs/_2371_ ),
    .Y(\soc/cpu/cpuregs/_2417_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4234_  (.A0(\soc/cpu/cpuregs/regs[26][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0256_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4235_  (.A0(\soc/cpu/cpuregs/regs[26][1] ),
    .A1(net130),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0257_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4236_  (.A0(\soc/cpu/cpuregs/regs[26][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0258_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4237_  (.A0(\soc/cpu/cpuregs/regs[26][3] ),
    .A1(net129),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0259_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4238_  (.A0(\soc/cpu/cpuregs/regs[26][4] ),
    .A1(net128),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0260_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4239_  (.A0(\soc/cpu/cpuregs/regs[26][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0261_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4240_  (.A0(\soc/cpu/cpuregs/regs[26][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0262_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4241_  (.A0(\soc/cpu/cpuregs/regs[26][7] ),
    .A1(net125),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0263_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4242_  (.A0(\soc/cpu/cpuregs/regs[26][8] ),
    .A1(net127),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0264_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4243_  (.A0(\soc/cpu/cpuregs/regs[26][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0265_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4245_  (.A0(\soc/cpu/cpuregs/regs[26][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0266_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4246_  (.A0(\soc/cpu/cpuregs/regs[26][11] ),
    .A1(net124),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0267_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4247_  (.A0(\soc/cpu/cpuregs/regs[26][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0268_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4248_  (.A0(\soc/cpu/cpuregs/regs[26][13] ),
    .A1(net105),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0269_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4249_  (.A0(\soc/cpu/cpuregs/regs[26][14] ),
    .A1(net114),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0270_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4250_  (.A0(\soc/cpu/cpuregs/regs[26][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0271_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4251_  (.A0(\soc/cpu/cpuregs/regs[26][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0272_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4252_  (.A0(\soc/cpu/cpuregs/regs[26][17] ),
    .A1(net88),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0273_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4253_  (.A0(\soc/cpu/cpuregs/regs[26][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0274_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4254_  (.A0(\soc/cpu/cpuregs/regs[26][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0275_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4256_  (.A0(\soc/cpu/cpuregs/regs[26][20] ),
    .A1(net64),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0276_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4257_  (.A0(\soc/cpu/cpuregs/regs[26][21] ),
    .A1(net59),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0277_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4258_  (.A0(\soc/cpu/cpuregs/regs[26][22] ),
    .A1(net60),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0278_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4259_  (.A0(\soc/cpu/cpuregs/regs[26][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0279_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4260_  (.A0(\soc/cpu/cpuregs/regs[26][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0280_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4261_  (.A0(\soc/cpu/cpuregs/regs[26][25] ),
    .A1(net58),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0281_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4262_  (.A0(\soc/cpu/cpuregs/regs[26][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0282_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4263_  (.A0(\soc/cpu/cpuregs/regs[26][27] ),
    .A1(net55),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0283_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4264_  (.A0(\soc/cpu/cpuregs/regs[26][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0284_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4265_  (.A0(\soc/cpu/cpuregs/regs[26][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(\soc/cpu/cpuregs/_2417_ ),
    .X(\soc/cpu/cpuregs/_0285_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4266_  (.A0(\soc/cpu/cpuregs/regs[26][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0286_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4267_  (.A0(\soc/cpu/cpuregs/regs[26][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net84),
    .X(\soc/cpu/cpuregs/_0287_ ));
 sky130_fd_sc_hd__or2_4 \soc/cpu/cpuregs/_4268_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/cpuregs/_2316_ ),
    .X(\soc/cpu/cpuregs/_2421_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4269_  (.A(\soc/cpu/cpuregs/_2421_ ),
    .B(\soc/cpu/cpuregs/_2372_ ),
    .Y(\soc/cpu/cpuregs/_2422_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4271_  (.A0(\soc/cpu/cpuregs/regs[21][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0288_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4272_  (.A0(\soc/cpu/cpuregs/regs[21][1] ),
    .A1(net130),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0289_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4273_  (.A0(\soc/cpu/cpuregs/regs[21][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0290_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4274_  (.A0(\soc/cpu/cpuregs/regs[21][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0291_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4275_  (.A0(\soc/cpu/cpuregs/regs[21][4] ),
    .A1(net128),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0292_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4276_  (.A0(\soc/cpu/cpuregs/regs[21][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0293_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4277_  (.A0(\soc/cpu/cpuregs/regs[21][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0294_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4278_  (.A0(\soc/cpu/cpuregs/regs[21][7] ),
    .A1(net125),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0295_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4279_  (.A0(\soc/cpu/cpuregs/regs[21][8] ),
    .A1(net126),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0296_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4280_  (.A0(\soc/cpu/cpuregs/regs[21][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0297_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4282_  (.A0(\soc/cpu/cpuregs/regs[21][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0298_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4283_  (.A0(\soc/cpu/cpuregs/regs[21][11] ),
    .A1(net123),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0299_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4284_  (.A0(\soc/cpu/cpuregs/regs[21][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0300_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4285_  (.A0(\soc/cpu/cpuregs/regs[21][13] ),
    .A1(net105),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0301_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4286_  (.A0(\soc/cpu/cpuregs/regs[21][14] ),
    .A1(net113),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0302_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4287_  (.A0(\soc/cpu/cpuregs/regs[21][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0303_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4288_  (.A0(\soc/cpu/cpuregs/regs[21][16] ),
    .A1(net69),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0304_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4289_  (.A0(\soc/cpu/cpuregs/regs[21][17] ),
    .A1(net87),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0305_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4290_  (.A0(\soc/cpu/cpuregs/regs[21][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0306_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4291_  (.A0(\soc/cpu/cpuregs/regs[21][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0307_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4293_  (.A0(\soc/cpu/cpuregs/regs[21][20] ),
    .A1(net64),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0308_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4294_  (.A0(\soc/cpu/cpuregs/regs[21][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0309_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4295_  (.A0(\soc/cpu/cpuregs/regs[21][22] ),
    .A1(net61),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0310_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4296_  (.A0(\soc/cpu/cpuregs/regs[21][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0311_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4297_  (.A0(\soc/cpu/cpuregs/regs[21][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0312_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4298_  (.A0(\soc/cpu/cpuregs/regs[21][25] ),
    .A1(net57),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0313_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4299_  (.A0(\soc/cpu/cpuregs/regs[21][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0314_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4300_  (.A0(\soc/cpu/cpuregs/regs[21][27] ),
    .A1(net55),
    .S(net82),
    .X(\soc/cpu/cpuregs/_0315_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4301_  (.A0(\soc/cpu/cpuregs/regs[21][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0316_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4302_  (.A0(\soc/cpu/cpuregs/regs[21][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0317_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4303_  (.A0(\soc/cpu/cpuregs/regs[21][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2422_ ),
    .X(\soc/cpu/cpuregs/_0318_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4304_  (.A0(\soc/cpu/cpuregs/regs[21][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net83),
    .X(\soc/cpu/cpuregs/_0319_ ));
 sky130_fd_sc_hd__nand3_4 \soc/cpu/cpuregs/_4305_  (.A(\soc/cpu/cpuregs_waddr[2] ),
    .B(\soc/cpu/cpuregs_waddr[3] ),
    .C(\soc/cpu/cpuregs_waddr[4] ),
    .Y(\soc/cpu/cpuregs/_2426_ ));
 sky130_fd_sc_hd__nor2_1 \soc/cpu/cpuregs/_4306_  (.A(\soc/cpu/cpuregs/_2371_ ),
    .B(\soc/cpu/cpuregs/_2426_ ),
    .Y(\soc/cpu/cpuregs/_2427_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4308_  (.A0(\soc/cpu/cpuregs/regs[30][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0320_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4309_  (.A0(\soc/cpu/cpuregs/regs[30][1] ),
    .A1(net130),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0321_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4310_  (.A0(\soc/cpu/cpuregs/regs[30][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0322_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4311_  (.A0(\soc/cpu/cpuregs/regs[30][3] ),
    .A1(net129),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0323_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4312_  (.A0(\soc/cpu/cpuregs/regs[30][4] ),
    .A1(net128),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0324_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4313_  (.A0(\soc/cpu/cpuregs/regs[30][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0325_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4314_  (.A0(\soc/cpu/cpuregs/regs[30][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0326_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4315_  (.A0(\soc/cpu/cpuregs/regs[30][7] ),
    .A1(net125),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0327_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4316_  (.A0(\soc/cpu/cpuregs/regs[30][8] ),
    .A1(net127),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0328_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4317_  (.A0(\soc/cpu/cpuregs/regs[30][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0329_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4319_  (.A0(\soc/cpu/cpuregs/regs[30][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0330_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4320_  (.A0(\soc/cpu/cpuregs/regs[30][11] ),
    .A1(net124),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0331_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4321_  (.A0(\soc/cpu/cpuregs/regs[30][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0332_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4322_  (.A0(\soc/cpu/cpuregs/regs[30][13] ),
    .A1(net105),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0333_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4323_  (.A0(\soc/cpu/cpuregs/regs[30][14] ),
    .A1(net114),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0334_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4324_  (.A0(\soc/cpu/cpuregs/regs[30][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0335_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4325_  (.A0(\soc/cpu/cpuregs/regs[30][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0336_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4326_  (.A0(\soc/cpu/cpuregs/regs[30][17] ),
    .A1(net88),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0337_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4327_  (.A0(\soc/cpu/cpuregs/regs[30][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0338_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4328_  (.A0(\soc/cpu/cpuregs/regs[30][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0339_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4330_  (.A0(\soc/cpu/cpuregs/regs[30][20] ),
    .A1(net63),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0340_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4331_  (.A0(\soc/cpu/cpuregs/regs[30][21] ),
    .A1(net59),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0341_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4332_  (.A0(\soc/cpu/cpuregs/regs[30][22] ),
    .A1(net60),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0342_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4333_  (.A0(\soc/cpu/cpuregs/regs[30][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0343_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4334_  (.A0(\soc/cpu/cpuregs/regs[30][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0344_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4335_  (.A0(\soc/cpu/cpuregs/regs[30][25] ),
    .A1(net58),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0345_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4336_  (.A0(\soc/cpu/cpuregs/regs[30][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net80),
    .X(\soc/cpu/cpuregs/_0346_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4337_  (.A0(\soc/cpu/cpuregs/regs[30][27] ),
    .A1(net55),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0347_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4338_  (.A0(\soc/cpu/cpuregs/regs[30][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0348_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4339_  (.A0(\soc/cpu/cpuregs/regs[30][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0349_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4340_  (.A0(\soc/cpu/cpuregs/regs[30][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0350_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4341_  (.A0(\soc/cpu/cpuregs/regs[30][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net81),
    .X(\soc/cpu/cpuregs/_0351_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4342_  (.A(\soc/cpu/cpuregs/_2354_ ),
    .B(\soc/cpu/cpuregs/_2366_ ),
    .Y(\soc/cpu/cpuregs/_2431_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4344_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[2][0] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0352_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4345_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[2][1] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0353_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4346_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[2][2] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0354_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4347_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[2][3] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0355_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4348_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[2][4] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0356_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4349_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[2][5] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0357_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4350_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[2][6] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0358_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4351_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[2][7] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0359_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4352_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[2][8] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0360_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4353_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[2][9] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0361_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4355_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[2][10] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0362_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4356_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[2][11] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0363_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4357_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[2][12] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0364_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4358_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[2][13] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0365_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4359_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[2][14] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0366_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4360_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[2][15] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0367_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4361_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[2][16] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0368_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4362_  (.A0(net88),
    .A1(\soc/cpu/cpuregs/regs[2][17] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0369_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4363_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[2][18] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0370_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4364_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[2][19] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0371_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4366_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[2][20] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0372_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4367_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[2][21] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0373_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4368_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[2][22] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0374_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4369_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[2][23] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0375_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4370_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[2][24] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0376_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4371_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[2][25] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0377_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4372_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[2][26] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0378_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4373_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[2][27] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0379_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4374_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[2][28] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0380_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4375_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[2][29] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0381_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4376_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[2][30] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0382_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4377_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[2][31] ),
    .S(\soc/cpu/cpuregs/_2431_ ),
    .X(\soc/cpu/cpuregs/_0383_ ));
 sky130_fd_sc_hd__nor3b_4 \soc/cpu/cpuregs/_4378_  (.A(\soc/cpu/cpuregs_waddr[2] ),
    .B(\soc/cpu/cpuregs_waddr[4] ),
    .C_N(\soc/cpu/cpuregs_waddr[3] ),
    .Y(\soc/cpu/cpuregs/_2435_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4379_  (.A(\soc/cpu/cpuregs/_2317_ ),
    .B(\soc/cpu/cpuregs/_2435_ ),
    .Y(\soc/cpu/cpuregs/_2436_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4381_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[9][0] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0384_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4382_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[9][1] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0385_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4383_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[9][2] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0386_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4384_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[9][3] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0387_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4385_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[9][4] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0388_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4386_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[9][5] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0389_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4387_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[9][6] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0390_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4388_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[9][7] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0391_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4389_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[9][8] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0392_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4390_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[9][9] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0393_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4392_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[9][10] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0394_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4393_  (.A0(net124),
    .A1(\soc/cpu/cpuregs/regs[9][11] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0395_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4394_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[9][12] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0396_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4395_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[9][13] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0397_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4396_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[9][14] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0398_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4397_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[9][15] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0399_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4398_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[9][16] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0400_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4399_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[9][17] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0401_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4400_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[9][18] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0402_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4401_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[9][19] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0403_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4403_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[9][20] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0404_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4404_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[9][21] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0405_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4405_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[9][22] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0406_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4406_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[9][23] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0407_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4407_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[9][24] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0408_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4408_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[9][25] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0409_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4409_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[9][26] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0410_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4410_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[9][27] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0411_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4411_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[9][28] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0412_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4412_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[9][29] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0413_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4413_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[9][30] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0414_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4414_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[9][31] ),
    .S(\soc/cpu/cpuregs/_2436_ ),
    .X(\soc/cpu/cpuregs/_0415_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4415_  (.A(\soc/cpu/cpuregs/_2277_ ),
    .B(\soc/cpu/cpuregs/_2361_ ),
    .Y(\soc/cpu/cpuregs/_2440_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4417_  (.A0(\soc/cpu/cpuregs/regs[24][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0416_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4418_  (.A0(\soc/cpu/cpuregs/regs[24][1] ),
    .A1(net130),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0417_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4419_  (.A0(\soc/cpu/cpuregs/regs[24][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0418_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4420_  (.A0(\soc/cpu/cpuregs/regs[24][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0419_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4421_  (.A0(\soc/cpu/cpuregs/regs[24][4] ),
    .A1(net128),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0420_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4422_  (.A0(\soc/cpu/cpuregs/regs[24][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0421_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4423_  (.A0(\soc/cpu/cpuregs/regs[24][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0422_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4424_  (.A0(\soc/cpu/cpuregs/regs[24][7] ),
    .A1(net125),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0423_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4425_  (.A0(\soc/cpu/cpuregs/regs[24][8] ),
    .A1(net126),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0424_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4426_  (.A0(\soc/cpu/cpuregs/regs[24][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0425_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4428_  (.A0(\soc/cpu/cpuregs/regs[24][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0426_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4429_  (.A0(\soc/cpu/cpuregs/regs[24][11] ),
    .A1(net123),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0427_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4430_  (.A0(\soc/cpu/cpuregs/regs[24][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0428_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4431_  (.A0(\soc/cpu/cpuregs/regs[24][13] ),
    .A1(net105),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0429_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4432_  (.A0(\soc/cpu/cpuregs/regs[24][14] ),
    .A1(net114),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0430_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4433_  (.A0(\soc/cpu/cpuregs/regs[24][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0431_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4434_  (.A0(\soc/cpu/cpuregs/regs[24][16] ),
    .A1(net69),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0432_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4435_  (.A0(\soc/cpu/cpuregs/regs[24][17] ),
    .A1(net87),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0433_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4436_  (.A0(\soc/cpu/cpuregs/regs[24][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0434_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4437_  (.A0(\soc/cpu/cpuregs/regs[24][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0435_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4439_  (.A0(\soc/cpu/cpuregs/regs[24][20] ),
    .A1(net63),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0436_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4440_  (.A0(\soc/cpu/cpuregs/regs[24][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0437_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4441_  (.A0(\soc/cpu/cpuregs/regs[24][22] ),
    .A1(net60),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0438_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4442_  (.A0(\soc/cpu/cpuregs/regs[24][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0439_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4443_  (.A0(\soc/cpu/cpuregs/regs[24][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0440_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4444_  (.A0(\soc/cpu/cpuregs/regs[24][25] ),
    .A1(net58),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0441_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4445_  (.A0(\soc/cpu/cpuregs/regs[24][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net95),
    .X(\soc/cpu/cpuregs/_0442_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4446_  (.A0(\soc/cpu/cpuregs/regs[24][27] ),
    .A1(net55),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0443_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4447_  (.A0(\soc/cpu/cpuregs/regs[24][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0444_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4448_  (.A0(\soc/cpu/cpuregs/regs[24][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(net96),
    .X(\soc/cpu/cpuregs/_0445_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4449_  (.A0(\soc/cpu/cpuregs/regs[24][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0446_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4450_  (.A0(\soc/cpu/cpuregs/regs[24][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(\soc/cpu/cpuregs/_2440_ ),
    .X(\soc/cpu/cpuregs/_0447_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4451_  (.A(\soc/cpu/cpuregs/_2361_ ),
    .B(\soc/cpu/cpuregs/_2426_ ),
    .Y(\soc/cpu/cpuregs/_2444_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4453_  (.A0(\soc/cpu/cpuregs/regs[28][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0448_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4454_  (.A0(\soc/cpu/cpuregs/regs[28][1] ),
    .A1(net130),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0449_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4455_  (.A0(\soc/cpu/cpuregs/regs[28][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0450_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4456_  (.A0(\soc/cpu/cpuregs/regs[28][3] ),
    .A1(net129),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0451_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4457_  (.A0(\soc/cpu/cpuregs/regs[28][4] ),
    .A1(net128),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0452_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4458_  (.A0(\soc/cpu/cpuregs/regs[28][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0453_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4459_  (.A0(\soc/cpu/cpuregs/regs[28][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0454_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4460_  (.A0(\soc/cpu/cpuregs/regs[28][7] ),
    .A1(net125),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0455_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4461_  (.A0(\soc/cpu/cpuregs/regs[28][8] ),
    .A1(net126),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0456_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4462_  (.A0(\soc/cpu/cpuregs/regs[28][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0457_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4464_  (.A0(\soc/cpu/cpuregs/regs[28][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0458_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4465_  (.A0(\soc/cpu/cpuregs/regs[28][11] ),
    .A1(net123),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0459_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4466_  (.A0(\soc/cpu/cpuregs/regs[28][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0460_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4467_  (.A0(\soc/cpu/cpuregs/regs[28][13] ),
    .A1(net105),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0461_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4468_  (.A0(\soc/cpu/cpuregs/regs[28][14] ),
    .A1(net114),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0462_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4469_  (.A0(\soc/cpu/cpuregs/regs[28][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0463_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4470_  (.A0(\soc/cpu/cpuregs/regs[28][16] ),
    .A1(net69),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0464_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4471_  (.A0(\soc/cpu/cpuregs/regs[28][17] ),
    .A1(net87),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0465_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4472_  (.A0(\soc/cpu/cpuregs/regs[28][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0466_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4473_  (.A0(\soc/cpu/cpuregs/regs[28][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0467_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4475_  (.A0(\soc/cpu/cpuregs/regs[28][20] ),
    .A1(net63),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0468_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4476_  (.A0(\soc/cpu/cpuregs/regs[28][21] ),
    .A1(net59),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0469_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4477_  (.A0(\soc/cpu/cpuregs/regs[28][22] ),
    .A1(net60),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0470_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4478_  (.A0(\soc/cpu/cpuregs/regs[28][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0471_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4479_  (.A0(\soc/cpu/cpuregs/regs[28][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0472_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4480_  (.A0(\soc/cpu/cpuregs/regs[28][25] ),
    .A1(net58),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0473_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4481_  (.A0(\soc/cpu/cpuregs/regs[28][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0474_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4482_  (.A0(\soc/cpu/cpuregs/regs[28][27] ),
    .A1(net55),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0475_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4483_  (.A0(\soc/cpu/cpuregs/regs[28][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net93),
    .X(\soc/cpu/cpuregs/_0476_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4484_  (.A0(\soc/cpu/cpuregs/regs[28][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(\soc/cpu/cpuregs/_2444_ ),
    .X(\soc/cpu/cpuregs/_0477_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4485_  (.A0(\soc/cpu/cpuregs/regs[28][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0478_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4486_  (.A0(\soc/cpu/cpuregs/regs[28][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net94),
    .X(\soc/cpu/cpuregs/_0479_ ));
 sky130_fd_sc_hd__and2_4 \soc/cpu/cpuregs/_4487_  (.A(\soc/cpu/_00074_ ),
    .B(\soc/cpu/cpuregs/_2360_ ),
    .X(\soc/cpu/cpuregs/_2448_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4488_  (.A(\soc/cpu/cpuregs/_2448_ ),
    .B(\soc/cpu/cpuregs/_2435_ ),
    .Y(\soc/cpu/cpuregs/_2449_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4490_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[8][0] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0480_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4491_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[8][1] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0481_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4492_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[8][2] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0482_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4493_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[8][3] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0483_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4494_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[8][4] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0484_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4495_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[8][5] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0485_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4496_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[8][6] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0486_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4497_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[8][7] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0487_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4498_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[8][8] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0488_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4499_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[8][9] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0489_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4501_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[8][10] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0490_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4502_  (.A0(net124),
    .A1(\soc/cpu/cpuregs/regs[8][11] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0491_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4503_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[8][12] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0492_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4504_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[8][13] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0493_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4505_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[8][14] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0494_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4506_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[8][15] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0495_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4507_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[8][16] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0496_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4508_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[8][17] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0497_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4509_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[8][18] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0498_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4510_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[8][19] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0499_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4512_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[8][20] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0500_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4513_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[8][21] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0501_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4514_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[8][22] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0502_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4515_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[8][23] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0503_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4516_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[8][24] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0504_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4517_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[8][25] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0505_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4518_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[8][26] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0506_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4519_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[8][27] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0507_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4520_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[8][28] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0508_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4521_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[8][29] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0509_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4522_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[8][30] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0510_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4523_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[8][31] ),
    .S(\soc/cpu/cpuregs/_2449_ ),
    .X(\soc/cpu/cpuregs/_0511_ ));
 sky130_fd_sc_hd__and3_4 \soc/cpu/cpuregs/_4524_  (.A(\soc/cpu/cpuregs_waddr[1] ),
    .B(\soc/cpu/cpuregs_waddr[0] ),
    .C(\soc/cpu/_00074_ ),
    .X(\soc/cpu/cpuregs/_2453_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4525_  (.A(\soc/cpu/cpuregs/_2453_ ),
    .B(\soc/cpu/cpuregs/_2366_ ),
    .Y(\soc/cpu/cpuregs/_2454_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4527_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[3][0] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0512_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4528_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[3][1] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0513_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4529_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[3][2] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0514_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4530_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[3][3] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0515_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4531_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[3][4] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0516_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4532_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[3][5] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0517_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4533_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[3][6] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0518_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4534_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[3][7] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0519_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4535_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[3][8] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0520_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4536_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[3][9] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0521_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4538_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[3][10] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0522_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4539_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[3][11] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0523_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4540_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[3][12] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0524_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4541_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[3][13] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0525_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4542_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[3][14] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0526_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4543_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[3][15] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0527_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4544_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[3][16] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0528_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4545_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[3][17] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0529_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4546_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[3][18] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0530_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4547_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[3][19] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0531_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4549_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[3][20] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0532_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4550_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[3][21] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0533_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4551_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[3][22] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0534_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4552_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[3][23] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0535_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4553_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[3][24] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0536_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4554_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[3][25] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0537_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4555_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[3][26] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0538_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4556_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[3][27] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0539_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4557_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[3][28] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0540_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4558_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[3][29] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0541_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4559_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[3][30] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0542_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4560_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[3][31] ),
    .S(\soc/cpu/cpuregs/_2454_ ),
    .X(\soc/cpu/cpuregs/_0543_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4561_  (.A(\soc/cpu/cpuregs/_2448_ ),
    .B(\soc/cpu/cpuregs/_2366_ ),
    .Y(\soc/cpu/cpuregs/_2458_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4563_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[0][0] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0544_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4564_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[0][1] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0545_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4565_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[0][2] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0546_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4566_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[0][3] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0547_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4567_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[0][4] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0548_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4568_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[0][5] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0549_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4569_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[0][6] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0550_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4570_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[0][7] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0551_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4571_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[0][8] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0552_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4572_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[0][9] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0553_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4574_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[0][10] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0554_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4575_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[0][11] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0555_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4576_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[0][12] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0556_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4577_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[0][13] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0557_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4578_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[0][14] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0558_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4579_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[0][15] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0559_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4580_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[0][16] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0560_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4581_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[0][17] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0561_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4582_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[0][18] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0562_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4583_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[0][19] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0563_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4585_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[0][20] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0564_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4586_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[0][21] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0565_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4587_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[0][22] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0566_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4588_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[0][23] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0567_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4589_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[0][24] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0568_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4590_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[0][25] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0569_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4591_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[0][26] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0570_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4592_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[0][27] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0571_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4593_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[0][28] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0572_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4594_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[0][29] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0573_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4595_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[0][30] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0574_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4596_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[0][31] ),
    .S(\soc/cpu/cpuregs/_2458_ ),
    .X(\soc/cpu/cpuregs/_0575_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4597_  (.A(\soc/cpu/cpuregs/_2354_ ),
    .B(\soc/cpu/cpuregs/_2435_ ),
    .Y(\soc/cpu/cpuregs/_2462_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4599_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[10][0] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0576_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4600_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[10][1] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0577_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4601_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[10][2] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0578_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4602_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[10][3] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0579_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4603_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[10][4] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0580_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4604_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[10][5] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0581_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4605_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[10][6] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0582_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4606_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[10][7] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0583_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4607_  (.A0(net127),
    .A1(\soc/cpu/cpuregs/regs[10][8] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0584_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4608_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[10][9] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0585_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4610_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[10][10] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0586_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4611_  (.A0(net124),
    .A1(\soc/cpu/cpuregs/regs[10][11] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0587_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4612_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[10][12] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0588_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4613_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[10][13] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0589_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4614_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[10][14] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0590_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4615_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[10][15] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0591_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4616_  (.A0(\soc/cpu/cpuregs_wrdata[16] ),
    .A1(\soc/cpu/cpuregs/regs[10][16] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0592_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4617_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[10][17] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0593_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4618_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[10][18] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0594_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4619_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[10][19] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0595_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4621_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[10][20] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0596_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4622_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[10][21] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0597_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4623_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[10][22] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0598_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4624_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[10][23] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0599_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4625_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[10][24] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0600_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4626_  (.A0(net58),
    .A1(\soc/cpu/cpuregs/regs[10][25] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0601_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4627_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[10][26] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0602_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4628_  (.A0(net55),
    .A1(\soc/cpu/cpuregs/regs[10][27] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0603_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4629_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[10][28] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0604_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4630_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[10][29] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0605_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4631_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[10][30] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0606_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4632_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[10][31] ),
    .S(\soc/cpu/cpuregs/_2462_ ),
    .X(\soc/cpu/cpuregs/_0607_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4633_  (.A(\soc/cpu/cpuregs/_2421_ ),
    .B(\soc/cpu/cpuregs/_2359_ ),
    .Y(\soc/cpu/cpuregs/_2466_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4635_  (.A0(\soc/cpu/cpuregs/regs[13][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0608_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4636_  (.A0(\soc/cpu/cpuregs/regs[13][1] ),
    .A1(net130),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0609_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4637_  (.A0(\soc/cpu/cpuregs/regs[13][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0610_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4638_  (.A0(\soc/cpu/cpuregs/regs[13][3] ),
    .A1(net129),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0611_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4639_  (.A0(\soc/cpu/cpuregs/regs[13][4] ),
    .A1(net128),
    .S(\soc/cpu/cpuregs/_2466_ ),
    .X(\soc/cpu/cpuregs/_0612_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4640_  (.A0(\soc/cpu/cpuregs/regs[13][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(\soc/cpu/cpuregs/_2466_ ),
    .X(\soc/cpu/cpuregs/_0613_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4641_  (.A0(\soc/cpu/cpuregs/regs[13][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0614_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4642_  (.A0(\soc/cpu/cpuregs/regs[13][7] ),
    .A1(net125),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0615_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4643_  (.A0(\soc/cpu/cpuregs/regs[13][8] ),
    .A1(net126),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0616_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4644_  (.A0(\soc/cpu/cpuregs/regs[13][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0617_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4646_  (.A0(\soc/cpu/cpuregs/regs[13][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0618_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4647_  (.A0(\soc/cpu/cpuregs/regs[13][11] ),
    .A1(net124),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0619_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4648_  (.A0(\soc/cpu/cpuregs/regs[13][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0620_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4649_  (.A0(\soc/cpu/cpuregs/regs[13][13] ),
    .A1(net105),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0621_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4650_  (.A0(\soc/cpu/cpuregs/regs[13][14] ),
    .A1(net113),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0622_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4651_  (.A0(\soc/cpu/cpuregs/regs[13][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0623_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4652_  (.A0(\soc/cpu/cpuregs/regs[13][16] ),
    .A1(net69),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0624_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4653_  (.A0(\soc/cpu/cpuregs/regs[13][17] ),
    .A1(net87),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0625_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4654_  (.A0(\soc/cpu/cpuregs/regs[13][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0626_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4655_  (.A0(\soc/cpu/cpuregs/regs[13][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2466_ ),
    .X(\soc/cpu/cpuregs/_0627_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4657_  (.A0(\soc/cpu/cpuregs/regs[13][20] ),
    .A1(net63),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0628_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4658_  (.A0(\soc/cpu/cpuregs/regs[13][21] ),
    .A1(net59),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0629_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4659_  (.A0(\soc/cpu/cpuregs/regs[13][22] ),
    .A1(net61),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0630_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4660_  (.A0(\soc/cpu/cpuregs/regs[13][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(\soc/cpu/cpuregs/_2466_ ),
    .X(\soc/cpu/cpuregs/_0631_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4661_  (.A0(\soc/cpu/cpuregs/regs[13][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0632_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4662_  (.A0(\soc/cpu/cpuregs/regs[13][25] ),
    .A1(net57),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0633_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4663_  (.A0(\soc/cpu/cpuregs/regs[13][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0634_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4664_  (.A0(\soc/cpu/cpuregs/regs[13][27] ),
    .A1(net56),
    .S(\soc/cpu/cpuregs/_2466_ ),
    .X(\soc/cpu/cpuregs/_0635_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4665_  (.A0(\soc/cpu/cpuregs/regs[13][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net78),
    .X(\soc/cpu/cpuregs/_0636_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4666_  (.A0(\soc/cpu/cpuregs/regs[13][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2466_ ),
    .X(\soc/cpu/cpuregs/_0637_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4667_  (.A0(\soc/cpu/cpuregs/regs[13][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0638_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4668_  (.A0(\soc/cpu/cpuregs/regs[13][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net79),
    .X(\soc/cpu/cpuregs/_0639_ ));
 sky130_fd_sc_hd__nor2_4 \soc/cpu/cpuregs/_4669_  (.A(\soc/cpu/cpuregs/_2277_ ),
    .B(\soc/cpu/cpuregs/_2421_ ),
    .Y(\soc/cpu/cpuregs/_2470_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4671_  (.A0(\soc/cpu/cpuregs/regs[25][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0640_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4672_  (.A0(\soc/cpu/cpuregs/regs[25][1] ),
    .A1(net130),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0641_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4673_  (.A0(\soc/cpu/cpuregs/regs[25][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0642_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4674_  (.A0(\soc/cpu/cpuregs/regs[25][3] ),
    .A1(net129),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0643_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4675_  (.A0(\soc/cpu/cpuregs/regs[25][4] ),
    .A1(net128),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0644_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4676_  (.A0(\soc/cpu/cpuregs/regs[25][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0645_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4677_  (.A0(\soc/cpu/cpuregs/regs[25][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0646_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4678_  (.A0(\soc/cpu/cpuregs/regs[25][7] ),
    .A1(net125),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0647_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4679_  (.A0(\soc/cpu/cpuregs/regs[25][8] ),
    .A1(net126),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0648_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4680_  (.A0(\soc/cpu/cpuregs/regs[25][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0649_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4682_  (.A0(\soc/cpu/cpuregs/regs[25][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0650_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4683_  (.A0(\soc/cpu/cpuregs/regs[25][11] ),
    .A1(net123),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0651_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4684_  (.A0(\soc/cpu/cpuregs/regs[25][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0652_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4685_  (.A0(\soc/cpu/cpuregs/regs[25][13] ),
    .A1(net105),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0653_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4686_  (.A0(\soc/cpu/cpuregs/regs[25][14] ),
    .A1(net114),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0654_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4687_  (.A0(\soc/cpu/cpuregs/regs[25][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0655_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4688_  (.A0(\soc/cpu/cpuregs/regs[25][16] ),
    .A1(net69),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0656_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4689_  (.A0(\soc/cpu/cpuregs/regs[25][17] ),
    .A1(net87),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0657_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4690_  (.A0(\soc/cpu/cpuregs/regs[25][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0658_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4691_  (.A0(\soc/cpu/cpuregs/regs[25][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0659_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4693_  (.A0(\soc/cpu/cpuregs/regs[25][20] ),
    .A1(net63),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0660_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4694_  (.A0(\soc/cpu/cpuregs/regs[25][21] ),
    .A1(net59),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0661_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4695_  (.A0(\soc/cpu/cpuregs/regs[25][22] ),
    .A1(net60),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0662_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4696_  (.A0(\soc/cpu/cpuregs/regs[25][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0663_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4697_  (.A0(\soc/cpu/cpuregs/regs[25][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0664_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4698_  (.A0(\soc/cpu/cpuregs/regs[25][25] ),
    .A1(net58),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0665_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4699_  (.A0(\soc/cpu/cpuregs/regs[25][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0666_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4700_  (.A0(\soc/cpu/cpuregs/regs[25][27] ),
    .A1(net55),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0667_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4701_  (.A0(\soc/cpu/cpuregs/regs[25][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net76),
    .X(\soc/cpu/cpuregs/_0668_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4702_  (.A0(\soc/cpu/cpuregs/regs[25][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(\soc/cpu/cpuregs/_2470_ ),
    .X(\soc/cpu/cpuregs/_0669_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4703_  (.A0(\soc/cpu/cpuregs/regs[25][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0670_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4704_  (.A0(\soc/cpu/cpuregs/regs[25][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net77),
    .X(\soc/cpu/cpuregs/_0671_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4705_  (.A(\soc/cpu/cpuregs/_2278_ ),
    .B(\soc/cpu/cpuregs/_2426_ ),
    .Y(\soc/cpu/cpuregs/_2474_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4707_  (.A0(\soc/cpu/cpuregs/regs[31][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0672_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4708_  (.A0(\soc/cpu/cpuregs/regs[31][1] ),
    .A1(net130),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0673_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4709_  (.A0(\soc/cpu/cpuregs/regs[31][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0674_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4710_  (.A0(\soc/cpu/cpuregs/regs[31][3] ),
    .A1(net129),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0675_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4711_  (.A0(\soc/cpu/cpuregs/regs[31][4] ),
    .A1(net128),
    .S(\soc/cpu/cpuregs/_2474_ ),
    .X(\soc/cpu/cpuregs/_0676_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4712_  (.A0(\soc/cpu/cpuregs/regs[31][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(\soc/cpu/cpuregs/_2474_ ),
    .X(\soc/cpu/cpuregs/_0677_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4713_  (.A0(\soc/cpu/cpuregs/regs[31][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0678_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4714_  (.A0(\soc/cpu/cpuregs/regs[31][7] ),
    .A1(net125),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0679_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4715_  (.A0(\soc/cpu/cpuregs/regs[31][8] ),
    .A1(net127),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0680_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4716_  (.A0(\soc/cpu/cpuregs/regs[31][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0681_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4718_  (.A0(\soc/cpu/cpuregs/regs[31][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0682_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4719_  (.A0(\soc/cpu/cpuregs/regs[31][11] ),
    .A1(net124),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0683_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4720_  (.A0(\soc/cpu/cpuregs/regs[31][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0684_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4721_  (.A0(\soc/cpu/cpuregs/regs[31][13] ),
    .A1(net105),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0685_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4722_  (.A0(\soc/cpu/cpuregs/regs[31][14] ),
    .A1(net114),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0686_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4723_  (.A0(\soc/cpu/cpuregs/regs[31][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0687_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4724_  (.A0(\soc/cpu/cpuregs/regs[31][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0688_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4725_  (.A0(\soc/cpu/cpuregs/regs[31][17] ),
    .A1(net88),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0689_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4726_  (.A0(\soc/cpu/cpuregs/regs[31][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0690_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4727_  (.A0(\soc/cpu/cpuregs/regs[31][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0691_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4729_  (.A0(\soc/cpu/cpuregs/regs[31][20] ),
    .A1(net63),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0692_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4730_  (.A0(\soc/cpu/cpuregs/regs[31][21] ),
    .A1(net59),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0693_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4731_  (.A0(\soc/cpu/cpuregs/regs[31][22] ),
    .A1(net60),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0694_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4732_  (.A0(\soc/cpu/cpuregs/regs[31][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(\soc/cpu/cpuregs/_2474_ ),
    .X(\soc/cpu/cpuregs/_0695_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4733_  (.A0(\soc/cpu/cpuregs/regs[31][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0696_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4734_  (.A0(\soc/cpu/cpuregs/regs[31][25] ),
    .A1(net58),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0697_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4735_  (.A0(\soc/cpu/cpuregs/regs[31][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net91),
    .X(\soc/cpu/cpuregs/_0698_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4736_  (.A0(\soc/cpu/cpuregs/regs[31][27] ),
    .A1(net55),
    .S(\soc/cpu/cpuregs/_2474_ ),
    .X(\soc/cpu/cpuregs/_0699_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4737_  (.A0(\soc/cpu/cpuregs/regs[31][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(\soc/cpu/cpuregs/_2474_ ),
    .X(\soc/cpu/cpuregs/_0700_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4738_  (.A0(\soc/cpu/cpuregs/regs[31][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0701_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4739_  (.A0(\soc/cpu/cpuregs/regs[31][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0702_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4740_  (.A0(\soc/cpu/cpuregs/regs[31][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net92),
    .X(\soc/cpu/cpuregs/_0703_ ));
 sky130_fd_sc_hd__nor3b_4 \soc/cpu/cpuregs/_4741_  (.A(\soc/cpu/cpuregs_waddr[2] ),
    .B(\soc/cpu/cpuregs_waddr[3] ),
    .C_N(\soc/cpu/cpuregs_waddr[4] ),
    .Y(\soc/cpu/cpuregs/_2478_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4742_  (.A(\soc/cpu/cpuregs/_2453_ ),
    .B(\soc/cpu/cpuregs/_2478_ ),
    .Y(\soc/cpu/cpuregs/_2479_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4744_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[19][0] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0704_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4745_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[19][1] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0705_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4746_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[19][2] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0706_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4747_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[19][3] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0707_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4748_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[19][4] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0708_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4749_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[19][5] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0709_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4750_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[19][6] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0710_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4751_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[19][7] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0711_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4752_  (.A0(net127),
    .A1(\soc/cpu/cpuregs/regs[19][8] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0712_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4753_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[19][9] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0713_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4755_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[19][10] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0714_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4756_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[19][11] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0715_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4757_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[19][12] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0716_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4758_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[19][13] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0717_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4759_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[19][14] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0718_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4760_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[19][15] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0719_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4761_  (.A0(\soc/cpu/cpuregs_wrdata[16] ),
    .A1(\soc/cpu/cpuregs/regs[19][16] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0720_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4762_  (.A0(net88),
    .A1(\soc/cpu/cpuregs/regs[19][17] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0721_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4763_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[19][18] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0722_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4764_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[19][19] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0723_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4766_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[19][20] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0724_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4767_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[19][21] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0725_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4768_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[19][22] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0726_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4769_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[19][23] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0727_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4770_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[19][24] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0728_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4771_  (.A0(net58),
    .A1(\soc/cpu/cpuregs/regs[19][25] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0729_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4772_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[19][26] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0730_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4773_  (.A0(net55),
    .A1(\soc/cpu/cpuregs/regs[19][27] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0731_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4774_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[19][28] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0732_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4775_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[19][29] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0733_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4776_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[19][30] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0734_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4777_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[19][31] ),
    .S(\soc/cpu/cpuregs/_2479_ ),
    .X(\soc/cpu/cpuregs/_0735_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4778_  (.A(\soc/cpu/cpuregs/_2453_ ),
    .B(\soc/cpu/cpuregs/_2435_ ),
    .Y(\soc/cpu/cpuregs/_2483_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4780_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[11][0] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0736_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4781_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[11][1] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0737_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4782_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[11][2] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0738_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4783_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[11][3] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0739_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4784_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[11][4] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0740_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4785_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[11][5] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0741_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4786_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[11][6] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0742_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4787_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[11][7] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0743_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4788_  (.A0(net127),
    .A1(\soc/cpu/cpuregs/regs[11][8] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0744_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4789_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[11][9] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0745_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4791_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[11][10] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0746_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4792_  (.A0(net124),
    .A1(\soc/cpu/cpuregs/regs[11][11] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0747_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4793_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[11][12] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0748_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4794_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[11][13] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0749_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4795_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[11][14] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0750_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4796_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[11][15] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0751_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4797_  (.A0(\soc/cpu/cpuregs_wrdata[16] ),
    .A1(\soc/cpu/cpuregs/regs[11][16] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0752_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4798_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[11][17] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0753_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4799_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[11][18] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0754_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4800_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[11][19] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0755_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4802_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[11][20] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0756_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4803_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[11][21] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0757_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4804_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[11][22] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0758_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4805_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[11][23] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0759_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4806_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[11][24] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0760_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4807_  (.A0(net58),
    .A1(\soc/cpu/cpuregs/regs[11][25] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0761_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4808_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[11][26] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0762_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4809_  (.A0(net55),
    .A1(\soc/cpu/cpuregs/regs[11][27] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0763_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4810_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[11][28] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0764_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4811_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[11][29] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0765_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4812_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[11][30] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0766_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4813_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[11][31] ),
    .S(\soc/cpu/cpuregs/_2483_ ),
    .X(\soc/cpu/cpuregs/_0767_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4814_  (.A(\soc/cpu/cpuregs/_2371_ ),
    .B(\soc/cpu/cpuregs/_2359_ ),
    .Y(\soc/cpu/cpuregs/_2487_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4816_  (.A0(\soc/cpu/cpuregs/regs[14][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0768_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4817_  (.A0(\soc/cpu/cpuregs/regs[14][1] ),
    .A1(net130),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0769_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4818_  (.A0(\soc/cpu/cpuregs/regs[14][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0770_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4819_  (.A0(\soc/cpu/cpuregs/regs[14][3] ),
    .A1(net129),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0771_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4820_  (.A0(\soc/cpu/cpuregs/regs[14][4] ),
    .A1(net128),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0772_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4821_  (.A0(\soc/cpu/cpuregs/regs[14][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0773_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4822_  (.A0(\soc/cpu/cpuregs/regs[14][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0774_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4823_  (.A0(\soc/cpu/cpuregs/regs[14][7] ),
    .A1(net125),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0775_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4824_  (.A0(\soc/cpu/cpuregs/regs[14][8] ),
    .A1(net127),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0776_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4825_  (.A0(\soc/cpu/cpuregs/regs[14][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0777_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4827_  (.A0(\soc/cpu/cpuregs/regs[14][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0778_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4828_  (.A0(\soc/cpu/cpuregs/regs[14][11] ),
    .A1(net124),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0779_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4829_  (.A0(\soc/cpu/cpuregs/regs[14][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0780_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4830_  (.A0(\soc/cpu/cpuregs/regs[14][13] ),
    .A1(net105),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0781_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4831_  (.A0(\soc/cpu/cpuregs/regs[14][14] ),
    .A1(net113),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0782_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4832_  (.A0(\soc/cpu/cpuregs/regs[14][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0783_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4833_  (.A0(\soc/cpu/cpuregs/regs[14][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0784_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4834_  (.A0(\soc/cpu/cpuregs/regs[14][17] ),
    .A1(net87),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0785_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4835_  (.A0(\soc/cpu/cpuregs/regs[14][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0786_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4836_  (.A0(\soc/cpu/cpuregs/regs[14][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0787_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4838_  (.A0(\soc/cpu/cpuregs/regs[14][20] ),
    .A1(net63),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0788_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4839_  (.A0(\soc/cpu/cpuregs/regs[14][21] ),
    .A1(net59),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0789_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4840_  (.A0(\soc/cpu/cpuregs/regs[14][22] ),
    .A1(net61),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0790_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4841_  (.A0(\soc/cpu/cpuregs/regs[14][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0791_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4842_  (.A0(\soc/cpu/cpuregs/regs[14][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0792_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4843_  (.A0(\soc/cpu/cpuregs/regs[14][25] ),
    .A1(net58),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0793_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4844_  (.A0(\soc/cpu/cpuregs/regs[14][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0794_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4845_  (.A0(\soc/cpu/cpuregs/regs[14][27] ),
    .A1(net55),
    .S(net74),
    .X(\soc/cpu/cpuregs/_0795_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4846_  (.A0(\soc/cpu/cpuregs/regs[14][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0796_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4847_  (.A0(\soc/cpu/cpuregs/regs[14][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(net75),
    .X(\soc/cpu/cpuregs/_0797_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4848_  (.A0(\soc/cpu/cpuregs/regs[14][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0798_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4849_  (.A0(\soc/cpu/cpuregs/regs[14][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(\soc/cpu/cpuregs/_2487_ ),
    .X(\soc/cpu/cpuregs/_0799_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4850_  (.A(\soc/cpu/cpuregs/_2315_ ),
    .B(\soc/cpu/cpuregs/_2448_ ),
    .Y(\soc/cpu/cpuregs/_2491_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4852_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[4][0] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0800_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4853_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[4][1] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0801_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4854_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[4][2] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0802_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4855_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[4][3] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0803_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4856_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[4][4] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0804_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4857_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[4][5] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0805_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4858_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[4][6] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0806_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4859_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[4][7] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0807_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4860_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[4][8] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0808_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4861_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[4][9] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0809_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4863_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[4][10] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0810_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4864_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[4][11] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0811_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4865_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[4][12] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0812_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4866_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[4][13] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0813_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4867_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[4][14] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0814_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4868_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[4][15] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0815_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4869_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[4][16] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0816_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4870_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[4][17] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0817_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4871_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[4][18] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0818_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4872_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[4][19] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0819_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4874_  (.A0(net63),
    .A1(\soc/cpu/cpuregs/regs[4][20] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0820_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4875_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[4][21] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0821_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4876_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[4][22] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0822_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4877_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[4][23] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0823_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4878_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[4][24] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0824_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4879_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[4][25] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0825_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4880_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[4][26] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0826_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4881_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[4][27] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0827_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4882_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[4][28] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0828_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4883_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[4][29] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0829_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4884_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[4][30] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0830_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4885_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[4][31] ),
    .S(\soc/cpu/cpuregs/_2491_ ),
    .X(\soc/cpu/cpuregs/_0831_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_4886_  (.A(\soc/cpu/cpuregs/_2278_ ),
    .B(\soc/cpu/cpuregs/_2359_ ),
    .Y(\soc/cpu/cpuregs/_2495_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4888_  (.A0(\soc/cpu/cpuregs/regs[15][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0832_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4889_  (.A0(\soc/cpu/cpuregs/regs[15][1] ),
    .A1(net130),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0833_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4890_  (.A0(\soc/cpu/cpuregs/regs[15][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0834_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4891_  (.A0(\soc/cpu/cpuregs/regs[15][3] ),
    .A1(net129),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0835_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4892_  (.A0(\soc/cpu/cpuregs/regs[15][4] ),
    .A1(net128),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0836_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4893_  (.A0(\soc/cpu/cpuregs/regs[15][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0837_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4894_  (.A0(\soc/cpu/cpuregs/regs[15][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0838_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4895_  (.A0(\soc/cpu/cpuregs/regs[15][7] ),
    .A1(net125),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0839_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4896_  (.A0(\soc/cpu/cpuregs/regs[15][8] ),
    .A1(net127),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0840_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4897_  (.A0(\soc/cpu/cpuregs/regs[15][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0841_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4899_  (.A0(\soc/cpu/cpuregs/regs[15][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0842_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4900_  (.A0(\soc/cpu/cpuregs/regs[15][11] ),
    .A1(net124),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0843_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4901_  (.A0(\soc/cpu/cpuregs/regs[15][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0844_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4902_  (.A0(\soc/cpu/cpuregs/regs[15][13] ),
    .A1(net105),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0845_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4903_  (.A0(\soc/cpu/cpuregs/regs[15][14] ),
    .A1(net113),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0846_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4904_  (.A0(\soc/cpu/cpuregs/regs[15][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0847_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4905_  (.A0(\soc/cpu/cpuregs/regs[15][16] ),
    .A1(\soc/cpu/cpuregs_wrdata[16] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0848_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4906_  (.A0(\soc/cpu/cpuregs/regs[15][17] ),
    .A1(net87),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0849_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4907_  (.A0(\soc/cpu/cpuregs/regs[15][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0850_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4908_  (.A0(\soc/cpu/cpuregs/regs[15][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0851_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4910_  (.A0(\soc/cpu/cpuregs/regs[15][20] ),
    .A1(net63),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0852_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4911_  (.A0(\soc/cpu/cpuregs/regs[15][21] ),
    .A1(net59),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0853_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4912_  (.A0(\soc/cpu/cpuregs/regs[15][22] ),
    .A1(net61),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0854_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4913_  (.A0(\soc/cpu/cpuregs/regs[15][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0855_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4914_  (.A0(\soc/cpu/cpuregs/regs[15][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0856_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4915_  (.A0(\soc/cpu/cpuregs/regs[15][25] ),
    .A1(net58),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0857_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4916_  (.A0(\soc/cpu/cpuregs/regs[15][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0858_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4917_  (.A0(\soc/cpu/cpuregs/regs[15][27] ),
    .A1(net55),
    .S(net89),
    .X(\soc/cpu/cpuregs/_0859_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4918_  (.A0(\soc/cpu/cpuregs/regs[15][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0860_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4919_  (.A0(\soc/cpu/cpuregs/regs[15][29] ),
    .A1(net52),
    .S(\soc/cpu/cpuregs/_2495_ ),
    .X(\soc/cpu/cpuregs/_0861_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4920_  (.A0(\soc/cpu/cpuregs/regs[15][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0862_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4921_  (.A0(\soc/cpu/cpuregs/regs[15][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net90),
    .X(\soc/cpu/cpuregs/_0863_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4922_  (.A(\soc/cpu/cpuregs/_2317_ ),
    .B(\soc/cpu/cpuregs/_2478_ ),
    .Y(\soc/cpu/cpuregs/_2499_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4924_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[17][0] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0864_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4925_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[17][1] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0865_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4926_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[17][2] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0866_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4927_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[17][3] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0867_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4928_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[17][4] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0868_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4929_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[17][5] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0869_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4930_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[17][6] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0870_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4931_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[17][7] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0871_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4932_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[17][8] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0872_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4933_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[17][9] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0873_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4935_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[17][10] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0874_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4936_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[17][11] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0875_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4937_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[17][12] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0876_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4938_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[17][13] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0877_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4939_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[17][14] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0878_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4940_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[17][15] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0879_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4941_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[17][16] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0880_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4942_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[17][17] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0881_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4943_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[17][18] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0882_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4944_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[17][19] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0883_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4946_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[17][20] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0884_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4947_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[17][21] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0885_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4948_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[17][22] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0886_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4949_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[17][23] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0887_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4950_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[17][24] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0888_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4951_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[17][25] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0889_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4952_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[17][26] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0890_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4953_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[17][27] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0891_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4954_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[17][28] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0892_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4955_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[17][29] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0893_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4956_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[17][30] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0894_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4957_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[17][31] ),
    .S(\soc/cpu/cpuregs/_2499_ ),
    .X(\soc/cpu/cpuregs/_0895_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4958_  (.A(\soc/cpu/cpuregs/_2354_ ),
    .B(\soc/cpu/cpuregs/_2478_ ),
    .Y(\soc/cpu/cpuregs/_2503_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4960_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[18][0] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0896_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4961_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[18][1] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0897_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4962_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[18][2] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0898_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4963_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[18][3] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0899_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4964_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[18][4] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0900_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4965_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[18][5] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0901_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4966_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[18][6] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0902_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4967_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[18][7] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0903_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4968_  (.A0(net127),
    .A1(\soc/cpu/cpuregs/regs[18][8] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0904_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4969_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[18][9] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0905_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4971_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[18][10] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0906_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4972_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[18][11] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0907_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4973_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[18][12] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0908_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4974_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[18][13] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0909_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4975_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[18][14] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0910_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4976_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[18][15] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0911_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4977_  (.A0(\soc/cpu/cpuregs_wrdata[16] ),
    .A1(\soc/cpu/cpuregs/regs[18][16] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0912_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4978_  (.A0(net88),
    .A1(\soc/cpu/cpuregs/regs[18][17] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0913_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4979_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[18][18] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0914_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4980_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[18][19] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0915_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4982_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[18][20] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0916_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4983_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[18][21] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0917_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4984_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[18][22] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0918_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4985_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[18][23] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0919_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4986_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[18][24] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0920_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4987_  (.A0(net58),
    .A1(\soc/cpu/cpuregs/regs[18][25] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0921_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4988_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[18][26] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0922_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4989_  (.A0(net55),
    .A1(\soc/cpu/cpuregs/regs[18][27] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0923_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4990_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[18][28] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0924_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4991_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[18][29] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0925_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4992_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[18][30] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0926_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4993_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[18][31] ),
    .S(\soc/cpu/cpuregs/_2503_ ),
    .X(\soc/cpu/cpuregs/_0927_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_4994_  (.A(\soc/cpu/cpuregs/_2453_ ),
    .B(\soc/cpu/cpuregs/_2315_ ),
    .Y(\soc/cpu/cpuregs/_2507_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4996_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[7][0] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0928_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4997_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[7][1] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0929_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4998_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[7][2] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0930_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_4999_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[7][3] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0931_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5000_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[7][4] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0932_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5001_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[7][5] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0933_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5002_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[7][6] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0934_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5003_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[7][7] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0935_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5004_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[7][8] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0936_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5005_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[7][9] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0937_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5007_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[7][10] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0938_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5008_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[7][11] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0939_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5009_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[7][12] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0940_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5010_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[7][13] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0941_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5011_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[7][14] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0942_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5012_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[7][15] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0943_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5013_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[7][16] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0944_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5014_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[7][17] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0945_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5015_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[7][18] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0946_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5016_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[7][19] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0947_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5018_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[7][20] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0948_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5019_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[7][21] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0949_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5020_  (.A0(net60),
    .A1(\soc/cpu/cpuregs/regs[7][22] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0950_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5021_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[7][23] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0951_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5022_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[7][24] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0952_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5023_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[7][25] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0953_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5024_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[7][26] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0954_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5025_  (.A0(net55),
    .A1(\soc/cpu/cpuregs/regs[7][27] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0955_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5026_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[7][28] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0956_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5027_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[7][29] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0957_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5028_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[7][30] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0958_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5029_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[7][31] ),
    .S(\soc/cpu/cpuregs/_2507_ ),
    .X(\soc/cpu/cpuregs/_0959_ ));
 sky130_fd_sc_hd__nor2_8 \soc/cpu/cpuregs/_5030_  (.A(\soc/cpu/cpuregs/_2421_ ),
    .B(\soc/cpu/cpuregs/_2426_ ),
    .Y(\soc/cpu/cpuregs/_2511_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5032_  (.A0(\soc/cpu/cpuregs/regs[29][0] ),
    .A1(\soc/cpu/cpuregs_wrdata[0] ),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0960_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5033_  (.A0(\soc/cpu/cpuregs/regs[29][1] ),
    .A1(net130),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0961_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5034_  (.A0(\soc/cpu/cpuregs/regs[29][2] ),
    .A1(\soc/cpu/cpuregs_wrdata[2] ),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0962_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5035_  (.A0(\soc/cpu/cpuregs/regs[29][3] ),
    .A1(net129),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0963_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5036_  (.A0(\soc/cpu/cpuregs/regs[29][4] ),
    .A1(net128),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0964_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5037_  (.A0(\soc/cpu/cpuregs/regs[29][5] ),
    .A1(\soc/cpu/cpuregs_wrdata[5] ),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0965_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5038_  (.A0(\soc/cpu/cpuregs/regs[29][6] ),
    .A1(\soc/cpu/cpuregs_wrdata[6] ),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0966_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5039_  (.A0(\soc/cpu/cpuregs/regs[29][7] ),
    .A1(net125),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0967_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5040_  (.A0(\soc/cpu/cpuregs/regs[29][8] ),
    .A1(net126),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0968_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5041_  (.A0(\soc/cpu/cpuregs/regs[29][9] ),
    .A1(\soc/cpu/cpuregs_wrdata[9] ),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0969_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5043_  (.A0(\soc/cpu/cpuregs/regs[29][10] ),
    .A1(\soc/cpu/cpuregs_wrdata[10] ),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0970_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5044_  (.A0(\soc/cpu/cpuregs/regs[29][11] ),
    .A1(net123),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0971_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5045_  (.A0(\soc/cpu/cpuregs/regs[29][12] ),
    .A1(\soc/cpu/cpuregs_wrdata[12] ),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0972_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5046_  (.A0(\soc/cpu/cpuregs/regs[29][13] ),
    .A1(net105),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0973_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5047_  (.A0(\soc/cpu/cpuregs/regs[29][14] ),
    .A1(net114),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0974_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5048_  (.A0(\soc/cpu/cpuregs/regs[29][15] ),
    .A1(\soc/cpu/cpuregs_wrdata[15] ),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0975_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5049_  (.A0(\soc/cpu/cpuregs/regs[29][16] ),
    .A1(net69),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0976_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5050_  (.A0(\soc/cpu/cpuregs/regs[29][17] ),
    .A1(net87),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0977_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5051_  (.A0(\soc/cpu/cpuregs/regs[29][18] ),
    .A1(\soc/cpu/cpuregs_wrdata[18] ),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0978_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5052_  (.A0(\soc/cpu/cpuregs/regs[29][19] ),
    .A1(\soc/cpu/cpuregs_wrdata[19] ),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0979_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5054_  (.A0(\soc/cpu/cpuregs/regs[29][20] ),
    .A1(net63),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0980_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5055_  (.A0(\soc/cpu/cpuregs/regs[29][21] ),
    .A1(net59),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0981_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5056_  (.A0(\soc/cpu/cpuregs/regs[29][22] ),
    .A1(net60),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0982_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5057_  (.A0(\soc/cpu/cpuregs/regs[29][23] ),
    .A1(\soc/cpu/cpuregs_wrdata[23] ),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0983_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5058_  (.A0(\soc/cpu/cpuregs/regs[29][24] ),
    .A1(\soc/cpu/cpuregs_wrdata[24] ),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0984_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5059_  (.A0(\soc/cpu/cpuregs/regs[29][25] ),
    .A1(net58),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0985_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5060_  (.A0(\soc/cpu/cpuregs/regs[29][26] ),
    .A1(\soc/cpu/cpuregs_wrdata[26] ),
    .S(net72),
    .X(\soc/cpu/cpuregs/_0986_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5061_  (.A0(\soc/cpu/cpuregs/regs[29][27] ),
    .A1(net55),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0987_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5062_  (.A0(\soc/cpu/cpuregs/regs[29][28] ),
    .A1(\soc/cpu/cpuregs_wrdata[28] ),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0988_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5063_  (.A0(\soc/cpu/cpuregs/regs[29][29] ),
    .A1(\soc/cpu/cpuregs_wrdata[29] ),
    .S(\soc/cpu/cpuregs/_2511_ ),
    .X(\soc/cpu/cpuregs/_0989_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5064_  (.A0(\soc/cpu/cpuregs/regs[29][30] ),
    .A1(\soc/cpu/cpuregs_wrdata[30] ),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0990_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5065_  (.A0(\soc/cpu/cpuregs/regs[29][31] ),
    .A1(\soc/cpu/cpuregs_wrdata[31] ),
    .S(net73),
    .X(\soc/cpu/cpuregs/_0991_ ));
 sky130_fd_sc_hd__nand2_8 \soc/cpu/cpuregs/_5066_  (.A(\soc/cpu/cpuregs/_2448_ ),
    .B(\soc/cpu/cpuregs/_2478_ ),
    .Y(\soc/cpu/cpuregs/_2515_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5068_  (.A0(\soc/cpu/cpuregs_wrdata[0] ),
    .A1(\soc/cpu/cpuregs/regs[16][0] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0992_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5069_  (.A0(net130),
    .A1(\soc/cpu/cpuregs/regs[16][1] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0993_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5070_  (.A0(\soc/cpu/cpuregs_wrdata[2] ),
    .A1(\soc/cpu/cpuregs/regs[16][2] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0994_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5071_  (.A0(net129),
    .A1(\soc/cpu/cpuregs/regs[16][3] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0995_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5072_  (.A0(net128),
    .A1(\soc/cpu/cpuregs/regs[16][4] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0996_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5073_  (.A0(\soc/cpu/cpuregs_wrdata[5] ),
    .A1(\soc/cpu/cpuregs/regs[16][5] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0997_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5074_  (.A0(\soc/cpu/cpuregs_wrdata[6] ),
    .A1(\soc/cpu/cpuregs/regs[16][6] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0998_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5075_  (.A0(net125),
    .A1(\soc/cpu/cpuregs/regs[16][7] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_0999_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5076_  (.A0(net126),
    .A1(\soc/cpu/cpuregs/regs[16][8] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1000_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5077_  (.A0(\soc/cpu/cpuregs_wrdata[9] ),
    .A1(\soc/cpu/cpuregs/regs[16][9] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1001_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5079_  (.A0(\soc/cpu/cpuregs_wrdata[10] ),
    .A1(\soc/cpu/cpuregs/regs[16][10] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1002_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5080_  (.A0(net123),
    .A1(\soc/cpu/cpuregs/regs[16][11] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1003_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5081_  (.A0(\soc/cpu/cpuregs_wrdata[12] ),
    .A1(\soc/cpu/cpuregs/regs[16][12] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1004_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5082_  (.A0(net105),
    .A1(\soc/cpu/cpuregs/regs[16][13] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1005_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5083_  (.A0(net113),
    .A1(\soc/cpu/cpuregs/regs[16][14] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1006_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5084_  (.A0(\soc/cpu/cpuregs_wrdata[15] ),
    .A1(\soc/cpu/cpuregs/regs[16][15] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1007_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5085_  (.A0(net69),
    .A1(\soc/cpu/cpuregs/regs[16][16] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1008_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5086_  (.A0(net87),
    .A1(\soc/cpu/cpuregs/regs[16][17] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1009_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5087_  (.A0(\soc/cpu/cpuregs_wrdata[18] ),
    .A1(\soc/cpu/cpuregs/regs[16][18] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1010_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5088_  (.A0(\soc/cpu/cpuregs_wrdata[19] ),
    .A1(\soc/cpu/cpuregs/regs[16][19] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1011_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5090_  (.A0(net64),
    .A1(\soc/cpu/cpuregs/regs[16][20] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1012_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5091_  (.A0(net59),
    .A1(\soc/cpu/cpuregs/regs[16][21] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1013_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5092_  (.A0(net61),
    .A1(\soc/cpu/cpuregs/regs[16][22] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1014_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5093_  (.A0(\soc/cpu/cpuregs_wrdata[23] ),
    .A1(\soc/cpu/cpuregs/regs[16][23] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1015_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5094_  (.A0(\soc/cpu/cpuregs_wrdata[24] ),
    .A1(\soc/cpu/cpuregs/regs[16][24] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1016_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5095_  (.A0(net57),
    .A1(\soc/cpu/cpuregs/regs[16][25] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1017_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5096_  (.A0(\soc/cpu/cpuregs_wrdata[26] ),
    .A1(\soc/cpu/cpuregs/regs[16][26] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1018_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5097_  (.A0(net56),
    .A1(\soc/cpu/cpuregs/regs[16][27] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1019_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5098_  (.A0(\soc/cpu/cpuregs_wrdata[28] ),
    .A1(\soc/cpu/cpuregs/regs[16][28] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1020_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5099_  (.A0(net52),
    .A1(\soc/cpu/cpuregs/regs[16][29] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1021_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5100_  (.A0(\soc/cpu/cpuregs_wrdata[30] ),
    .A1(\soc/cpu/cpuregs/regs[16][30] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1022_ ));
 sky130_fd_sc_hd__mux2_1 \soc/cpu/cpuregs/_5101_  (.A0(\soc/cpu/cpuregs_wrdata[31] ),
    .A1(\soc/cpu/cpuregs/regs[16][31] ),
    .S(\soc/cpu/cpuregs/_2515_ ),
    .X(\soc/cpu/cpuregs/_1023_ ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5102_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0000_ ),
    .Q(\soc/cpu/cpuregs/regs[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5103_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0001_ ),
    .Q(\soc/cpu/cpuregs/regs[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5104_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0002_ ),
    .Q(\soc/cpu/cpuregs/regs[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5105_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0003_ ),
    .Q(\soc/cpu/cpuregs/regs[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5106_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0004_ ),
    .Q(\soc/cpu/cpuregs/regs[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5107_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0005_ ),
    .Q(\soc/cpu/cpuregs/regs[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5108_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0006_ ),
    .Q(\soc/cpu/cpuregs/regs[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5109_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0007_ ),
    .Q(\soc/cpu/cpuregs/regs[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5110_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0008_ ),
    .Q(\soc/cpu/cpuregs/regs[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5111_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/cpuregs/_0009_ ),
    .Q(\soc/cpu/cpuregs/regs[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5112_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0010_ ),
    .Q(\soc/cpu/cpuregs/regs[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5113_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0011_ ),
    .Q(\soc/cpu/cpuregs/regs[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5114_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0012_ ),
    .Q(\soc/cpu/cpuregs/regs[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5115_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0013_ ),
    .Q(\soc/cpu/cpuregs/regs[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5116_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0014_ ),
    .Q(\soc/cpu/cpuregs/regs[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5117_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0015_ ),
    .Q(\soc/cpu/cpuregs/regs[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5118_  (.CLK(clknet_leaf_11_clk),
    .D(\soc/cpu/cpuregs/_0016_ ),
    .Q(\soc/cpu/cpuregs/regs[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5119_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0017_ ),
    .Q(\soc/cpu/cpuregs/regs[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5120_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0018_ ),
    .Q(\soc/cpu/cpuregs/regs[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5121_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0019_ ),
    .Q(\soc/cpu/cpuregs/regs[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5122_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0020_ ),
    .Q(\soc/cpu/cpuregs/regs[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5123_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0021_ ),
    .Q(\soc/cpu/cpuregs/regs[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5124_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0022_ ),
    .Q(\soc/cpu/cpuregs/regs[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5125_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0023_ ),
    .Q(\soc/cpu/cpuregs/regs[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5126_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0024_ ),
    .Q(\soc/cpu/cpuregs/regs[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5127_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0025_ ),
    .Q(\soc/cpu/cpuregs/regs[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5128_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0026_ ),
    .Q(\soc/cpu/cpuregs/regs[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5129_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0027_ ),
    .Q(\soc/cpu/cpuregs/regs[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5130_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0028_ ),
    .Q(\soc/cpu/cpuregs/regs[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5131_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0029_ ),
    .Q(\soc/cpu/cpuregs/regs[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5132_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0030_ ),
    .Q(\soc/cpu/cpuregs/regs[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5133_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0031_ ),
    .Q(\soc/cpu/cpuregs/regs[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5134_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0032_ ),
    .Q(\soc/cpu/cpuregs/regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5135_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0033_ ),
    .Q(\soc/cpu/cpuregs/regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5136_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0034_ ),
    .Q(\soc/cpu/cpuregs/regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5137_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0035_ ),
    .Q(\soc/cpu/cpuregs/regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5138_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0036_ ),
    .Q(\soc/cpu/cpuregs/regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5139_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0037_ ),
    .Q(\soc/cpu/cpuregs/regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5140_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0038_ ),
    .Q(\soc/cpu/cpuregs/regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5141_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0039_ ),
    .Q(\soc/cpu/cpuregs/regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5142_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0040_ ),
    .Q(\soc/cpu/cpuregs/regs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5143_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0041_ ),
    .Q(\soc/cpu/cpuregs/regs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5144_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0042_ ),
    .Q(\soc/cpu/cpuregs/regs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5145_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0043_ ),
    .Q(\soc/cpu/cpuregs/regs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5146_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0044_ ),
    .Q(\soc/cpu/cpuregs/regs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5147_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0045_ ),
    .Q(\soc/cpu/cpuregs/regs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5148_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0046_ ),
    .Q(\soc/cpu/cpuregs/regs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5149_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0047_ ),
    .Q(\soc/cpu/cpuregs/regs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5150_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0048_ ),
    .Q(\soc/cpu/cpuregs/regs[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5151_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0049_ ),
    .Q(\soc/cpu/cpuregs/regs[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5152_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0050_ ),
    .Q(\soc/cpu/cpuregs/regs[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5153_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0051_ ),
    .Q(\soc/cpu/cpuregs/regs[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5154_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0052_ ),
    .Q(\soc/cpu/cpuregs/regs[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5155_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0053_ ),
    .Q(\soc/cpu/cpuregs/regs[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5156_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0054_ ),
    .Q(\soc/cpu/cpuregs/regs[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5157_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0055_ ),
    .Q(\soc/cpu/cpuregs/regs[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5158_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0056_ ),
    .Q(\soc/cpu/cpuregs/regs[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5159_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0057_ ),
    .Q(\soc/cpu/cpuregs/regs[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5160_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0058_ ),
    .Q(\soc/cpu/cpuregs/regs[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5161_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0059_ ),
    .Q(\soc/cpu/cpuregs/regs[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5162_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0060_ ),
    .Q(\soc/cpu/cpuregs/regs[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5163_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0061_ ),
    .Q(\soc/cpu/cpuregs/regs[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5164_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0062_ ),
    .Q(\soc/cpu/cpuregs/regs[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5165_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0063_ ),
    .Q(\soc/cpu/cpuregs/regs[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5166_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0064_ ),
    .Q(\soc/cpu/cpuregs/regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5167_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0065_ ),
    .Q(\soc/cpu/cpuregs/regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5168_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0066_ ),
    .Q(\soc/cpu/cpuregs/regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5169_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0067_ ),
    .Q(\soc/cpu/cpuregs/regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5170_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0068_ ),
    .Q(\soc/cpu/cpuregs/regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5171_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0069_ ),
    .Q(\soc/cpu/cpuregs/regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5172_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0070_ ),
    .Q(\soc/cpu/cpuregs/regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5173_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0071_ ),
    .Q(\soc/cpu/cpuregs/regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5174_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0072_ ),
    .Q(\soc/cpu/cpuregs/regs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5175_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0073_ ),
    .Q(\soc/cpu/cpuregs/regs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5176_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0074_ ),
    .Q(\soc/cpu/cpuregs/regs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5177_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0075_ ),
    .Q(\soc/cpu/cpuregs/regs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5178_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0076_ ),
    .Q(\soc/cpu/cpuregs/regs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5179_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0077_ ),
    .Q(\soc/cpu/cpuregs/regs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5180_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0078_ ),
    .Q(\soc/cpu/cpuregs/regs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5181_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0079_ ),
    .Q(\soc/cpu/cpuregs/regs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5182_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0080_ ),
    .Q(\soc/cpu/cpuregs/regs[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5183_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0081_ ),
    .Q(\soc/cpu/cpuregs/regs[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5184_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0082_ ),
    .Q(\soc/cpu/cpuregs/regs[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5185_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0083_ ),
    .Q(\soc/cpu/cpuregs/regs[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5186_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0084_ ),
    .Q(\soc/cpu/cpuregs/regs[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5187_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0085_ ),
    .Q(\soc/cpu/cpuregs/regs[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5188_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0086_ ),
    .Q(\soc/cpu/cpuregs/regs[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5189_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0087_ ),
    .Q(\soc/cpu/cpuregs/regs[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5190_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0088_ ),
    .Q(\soc/cpu/cpuregs/regs[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5191_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0089_ ),
    .Q(\soc/cpu/cpuregs/regs[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5192_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0090_ ),
    .Q(\soc/cpu/cpuregs/regs[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5193_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0091_ ),
    .Q(\soc/cpu/cpuregs/regs[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5194_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0092_ ),
    .Q(\soc/cpu/cpuregs/regs[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5195_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0093_ ),
    .Q(\soc/cpu/cpuregs/regs[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5196_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0094_ ),
    .Q(\soc/cpu/cpuregs/regs[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5197_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0095_ ),
    .Q(\soc/cpu/cpuregs/regs[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5198_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0096_ ),
    .Q(\soc/cpu/cpuregs/regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5199_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0097_ ),
    .Q(\soc/cpu/cpuregs/regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5200_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0098_ ),
    .Q(\soc/cpu/cpuregs/regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5201_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0099_ ),
    .Q(\soc/cpu/cpuregs/regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5202_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0100_ ),
    .Q(\soc/cpu/cpuregs/regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5203_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0101_ ),
    .Q(\soc/cpu/cpuregs/regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5204_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0102_ ),
    .Q(\soc/cpu/cpuregs/regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5205_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0103_ ),
    .Q(\soc/cpu/cpuregs/regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5206_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0104_ ),
    .Q(\soc/cpu/cpuregs/regs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5207_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0105_ ),
    .Q(\soc/cpu/cpuregs/regs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5208_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0106_ ),
    .Q(\soc/cpu/cpuregs/regs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5209_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0107_ ),
    .Q(\soc/cpu/cpuregs/regs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5210_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0108_ ),
    .Q(\soc/cpu/cpuregs/regs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5211_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0109_ ),
    .Q(\soc/cpu/cpuregs/regs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5212_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0110_ ),
    .Q(\soc/cpu/cpuregs/regs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5213_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0111_ ),
    .Q(\soc/cpu/cpuregs/regs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5214_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0112_ ),
    .Q(\soc/cpu/cpuregs/regs[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5215_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0113_ ),
    .Q(\soc/cpu/cpuregs/regs[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5216_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0114_ ),
    .Q(\soc/cpu/cpuregs/regs[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5217_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0115_ ),
    .Q(\soc/cpu/cpuregs/regs[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5218_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0116_ ),
    .Q(\soc/cpu/cpuregs/regs[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5219_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0117_ ),
    .Q(\soc/cpu/cpuregs/regs[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5220_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0118_ ),
    .Q(\soc/cpu/cpuregs/regs[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5221_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0119_ ),
    .Q(\soc/cpu/cpuregs/regs[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5222_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0120_ ),
    .Q(\soc/cpu/cpuregs/regs[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5223_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0121_ ),
    .Q(\soc/cpu/cpuregs/regs[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5224_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0122_ ),
    .Q(\soc/cpu/cpuregs/regs[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5225_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0123_ ),
    .Q(\soc/cpu/cpuregs/regs[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5226_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0124_ ),
    .Q(\soc/cpu/cpuregs/regs[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5227_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0125_ ),
    .Q(\soc/cpu/cpuregs/regs[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5228_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0126_ ),
    .Q(\soc/cpu/cpuregs/regs[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5229_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0127_ ),
    .Q(\soc/cpu/cpuregs/regs[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5230_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0128_ ),
    .Q(\soc/cpu/cpuregs/regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5231_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0129_ ),
    .Q(\soc/cpu/cpuregs/regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5232_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0130_ ),
    .Q(\soc/cpu/cpuregs/regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5233_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0131_ ),
    .Q(\soc/cpu/cpuregs/regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5234_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0132_ ),
    .Q(\soc/cpu/cpuregs/regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5235_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0133_ ),
    .Q(\soc/cpu/cpuregs/regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5236_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0134_ ),
    .Q(\soc/cpu/cpuregs/regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5237_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0135_ ),
    .Q(\soc/cpu/cpuregs/regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5238_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0136_ ),
    .Q(\soc/cpu/cpuregs/regs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5239_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0137_ ),
    .Q(\soc/cpu/cpuregs/regs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5240_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0138_ ),
    .Q(\soc/cpu/cpuregs/regs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5241_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0139_ ),
    .Q(\soc/cpu/cpuregs/regs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5242_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0140_ ),
    .Q(\soc/cpu/cpuregs/regs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5243_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0141_ ),
    .Q(\soc/cpu/cpuregs/regs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5244_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0142_ ),
    .Q(\soc/cpu/cpuregs/regs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5245_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0143_ ),
    .Q(\soc/cpu/cpuregs/regs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5246_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0144_ ),
    .Q(\soc/cpu/cpuregs/regs[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5247_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0145_ ),
    .Q(\soc/cpu/cpuregs/regs[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5248_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0146_ ),
    .Q(\soc/cpu/cpuregs/regs[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5249_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0147_ ),
    .Q(\soc/cpu/cpuregs/regs[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5250_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0148_ ),
    .Q(\soc/cpu/cpuregs/regs[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5251_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0149_ ),
    .Q(\soc/cpu/cpuregs/regs[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5252_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0150_ ),
    .Q(\soc/cpu/cpuregs/regs[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5253_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0151_ ),
    .Q(\soc/cpu/cpuregs/regs[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5254_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0152_ ),
    .Q(\soc/cpu/cpuregs/regs[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5255_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0153_ ),
    .Q(\soc/cpu/cpuregs/regs[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5256_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0154_ ),
    .Q(\soc/cpu/cpuregs/regs[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5257_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0155_ ),
    .Q(\soc/cpu/cpuregs/regs[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5258_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0156_ ),
    .Q(\soc/cpu/cpuregs/regs[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5259_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0157_ ),
    .Q(\soc/cpu/cpuregs/regs[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5260_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0158_ ),
    .Q(\soc/cpu/cpuregs/regs[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5261_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0159_ ),
    .Q(\soc/cpu/cpuregs/regs[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5262_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0160_ ),
    .Q(\soc/cpu/cpuregs/regs[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5263_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0161_ ),
    .Q(\soc/cpu/cpuregs/regs[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5264_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0162_ ),
    .Q(\soc/cpu/cpuregs/regs[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5265_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0163_ ),
    .Q(\soc/cpu/cpuregs/regs[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5266_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0164_ ),
    .Q(\soc/cpu/cpuregs/regs[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5267_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0165_ ),
    .Q(\soc/cpu/cpuregs/regs[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5268_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0166_ ),
    .Q(\soc/cpu/cpuregs/regs[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5269_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0167_ ),
    .Q(\soc/cpu/cpuregs/regs[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5270_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0168_ ),
    .Q(\soc/cpu/cpuregs/regs[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5271_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/cpuregs/_0169_ ),
    .Q(\soc/cpu/cpuregs/regs[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5272_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0170_ ),
    .Q(\soc/cpu/cpuregs/regs[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5273_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0171_ ),
    .Q(\soc/cpu/cpuregs/regs[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5274_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0172_ ),
    .Q(\soc/cpu/cpuregs/regs[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5275_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0173_ ),
    .Q(\soc/cpu/cpuregs/regs[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5276_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0174_ ),
    .Q(\soc/cpu/cpuregs/regs[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5277_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0175_ ),
    .Q(\soc/cpu/cpuregs/regs[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5278_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0176_ ),
    .Q(\soc/cpu/cpuregs/regs[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5279_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0177_ ),
    .Q(\soc/cpu/cpuregs/regs[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5280_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0178_ ),
    .Q(\soc/cpu/cpuregs/regs[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5281_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0179_ ),
    .Q(\soc/cpu/cpuregs/regs[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5282_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0180_ ),
    .Q(\soc/cpu/cpuregs/regs[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5283_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0181_ ),
    .Q(\soc/cpu/cpuregs/regs[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5284_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0182_ ),
    .Q(\soc/cpu/cpuregs/regs[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5285_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0183_ ),
    .Q(\soc/cpu/cpuregs/regs[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5286_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0184_ ),
    .Q(\soc/cpu/cpuregs/regs[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5287_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0185_ ),
    .Q(\soc/cpu/cpuregs/regs[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5288_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0186_ ),
    .Q(\soc/cpu/cpuregs/regs[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5289_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0187_ ),
    .Q(\soc/cpu/cpuregs/regs[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5290_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0188_ ),
    .Q(\soc/cpu/cpuregs/regs[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5291_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0189_ ),
    .Q(\soc/cpu/cpuregs/regs[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5292_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0190_ ),
    .Q(\soc/cpu/cpuregs/regs[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5293_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0191_ ),
    .Q(\soc/cpu/cpuregs/regs[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5294_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0192_ ),
    .Q(\soc/cpu/cpuregs/regs[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5295_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0193_ ),
    .Q(\soc/cpu/cpuregs/regs[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5296_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0194_ ),
    .Q(\soc/cpu/cpuregs/regs[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5297_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0195_ ),
    .Q(\soc/cpu/cpuregs/regs[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5298_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0196_ ),
    .Q(\soc/cpu/cpuregs/regs[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5299_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0197_ ),
    .Q(\soc/cpu/cpuregs/regs[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5300_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0198_ ),
    .Q(\soc/cpu/cpuregs/regs[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5301_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0199_ ),
    .Q(\soc/cpu/cpuregs/regs[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5302_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0200_ ),
    .Q(\soc/cpu/cpuregs/regs[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5303_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/cpuregs/_0201_ ),
    .Q(\soc/cpu/cpuregs/regs[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5304_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0202_ ),
    .Q(\soc/cpu/cpuregs/regs[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5305_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0203_ ),
    .Q(\soc/cpu/cpuregs/regs[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5306_  (.CLK(clknet_leaf_11_clk),
    .D(\soc/cpu/cpuregs/_0204_ ),
    .Q(\soc/cpu/cpuregs/regs[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5307_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0205_ ),
    .Q(\soc/cpu/cpuregs/regs[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5308_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0206_ ),
    .Q(\soc/cpu/cpuregs/regs[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5309_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0207_ ),
    .Q(\soc/cpu/cpuregs/regs[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5310_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0208_ ),
    .Q(\soc/cpu/cpuregs/regs[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5311_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0209_ ),
    .Q(\soc/cpu/cpuregs/regs[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5312_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0210_ ),
    .Q(\soc/cpu/cpuregs/regs[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5313_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0211_ ),
    .Q(\soc/cpu/cpuregs/regs[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5314_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0212_ ),
    .Q(\soc/cpu/cpuregs/regs[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5315_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0213_ ),
    .Q(\soc/cpu/cpuregs/regs[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5316_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0214_ ),
    .Q(\soc/cpu/cpuregs/regs[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5317_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0215_ ),
    .Q(\soc/cpu/cpuregs/regs[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5318_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0216_ ),
    .Q(\soc/cpu/cpuregs/regs[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5319_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0217_ ),
    .Q(\soc/cpu/cpuregs/regs[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5320_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0218_ ),
    .Q(\soc/cpu/cpuregs/regs[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5321_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0219_ ),
    .Q(\soc/cpu/cpuregs/regs[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5322_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0220_ ),
    .Q(\soc/cpu/cpuregs/regs[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5323_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0221_ ),
    .Q(\soc/cpu/cpuregs/regs[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5324_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0222_ ),
    .Q(\soc/cpu/cpuregs/regs[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5325_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0223_ ),
    .Q(\soc/cpu/cpuregs/regs[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5326_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0224_ ),
    .Q(\soc/cpu/cpuregs/regs[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5327_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0225_ ),
    .Q(\soc/cpu/cpuregs/regs[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5328_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0226_ ),
    .Q(\soc/cpu/cpuregs/regs[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5329_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0227_ ),
    .Q(\soc/cpu/cpuregs/regs[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5330_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0228_ ),
    .Q(\soc/cpu/cpuregs/regs[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5331_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0229_ ),
    .Q(\soc/cpu/cpuregs/regs[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5332_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0230_ ),
    .Q(\soc/cpu/cpuregs/regs[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5333_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0231_ ),
    .Q(\soc/cpu/cpuregs/regs[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5334_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0232_ ),
    .Q(\soc/cpu/cpuregs/regs[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5335_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0233_ ),
    .Q(\soc/cpu/cpuregs/regs[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5336_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0234_ ),
    .Q(\soc/cpu/cpuregs/regs[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5337_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0235_ ),
    .Q(\soc/cpu/cpuregs/regs[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5338_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0236_ ),
    .Q(\soc/cpu/cpuregs/regs[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5339_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0237_ ),
    .Q(\soc/cpu/cpuregs/regs[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5340_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0238_ ),
    .Q(\soc/cpu/cpuregs/regs[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5341_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0239_ ),
    .Q(\soc/cpu/cpuregs/regs[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5342_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0240_ ),
    .Q(\soc/cpu/cpuregs/regs[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5343_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0241_ ),
    .Q(\soc/cpu/cpuregs/regs[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5344_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0242_ ),
    .Q(\soc/cpu/cpuregs/regs[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5345_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0243_ ),
    .Q(\soc/cpu/cpuregs/regs[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5346_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0244_ ),
    .Q(\soc/cpu/cpuregs/regs[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5347_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0245_ ),
    .Q(\soc/cpu/cpuregs/regs[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5348_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0246_ ),
    .Q(\soc/cpu/cpuregs/regs[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5349_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0247_ ),
    .Q(\soc/cpu/cpuregs/regs[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5350_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0248_ ),
    .Q(\soc/cpu/cpuregs/regs[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5351_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0249_ ),
    .Q(\soc/cpu/cpuregs/regs[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5352_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0250_ ),
    .Q(\soc/cpu/cpuregs/regs[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5353_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0251_ ),
    .Q(\soc/cpu/cpuregs/regs[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5354_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0252_ ),
    .Q(\soc/cpu/cpuregs/regs[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5355_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0253_ ),
    .Q(\soc/cpu/cpuregs/regs[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5356_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0254_ ),
    .Q(\soc/cpu/cpuregs/regs[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5357_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0255_ ),
    .Q(\soc/cpu/cpuregs/regs[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5358_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0256_ ),
    .Q(\soc/cpu/cpuregs/regs[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5359_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0257_ ),
    .Q(\soc/cpu/cpuregs/regs[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5360_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0258_ ),
    .Q(\soc/cpu/cpuregs/regs[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5361_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0259_ ),
    .Q(\soc/cpu/cpuregs/regs[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5362_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0260_ ),
    .Q(\soc/cpu/cpuregs/regs[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5363_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0261_ ),
    .Q(\soc/cpu/cpuregs/regs[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5364_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0262_ ),
    .Q(\soc/cpu/cpuregs/regs[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5365_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0263_ ),
    .Q(\soc/cpu/cpuregs/regs[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5366_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0264_ ),
    .Q(\soc/cpu/cpuregs/regs[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5367_  (.CLK(clknet_leaf_9_clk),
    .D(\soc/cpu/cpuregs/_0265_ ),
    .Q(\soc/cpu/cpuregs/regs[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5368_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0266_ ),
    .Q(\soc/cpu/cpuregs/regs[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5369_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0267_ ),
    .Q(\soc/cpu/cpuregs/regs[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5370_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0268_ ),
    .Q(\soc/cpu/cpuregs/regs[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5371_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0269_ ),
    .Q(\soc/cpu/cpuregs/regs[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5372_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0270_ ),
    .Q(\soc/cpu/cpuregs/regs[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5373_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0271_ ),
    .Q(\soc/cpu/cpuregs/regs[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5374_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0272_ ),
    .Q(\soc/cpu/cpuregs/regs[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5375_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0273_ ),
    .Q(\soc/cpu/cpuregs/regs[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5376_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0274_ ),
    .Q(\soc/cpu/cpuregs/regs[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5377_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0275_ ),
    .Q(\soc/cpu/cpuregs/regs[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5378_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0276_ ),
    .Q(\soc/cpu/cpuregs/regs[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5379_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0277_ ),
    .Q(\soc/cpu/cpuregs/regs[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5380_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0278_ ),
    .Q(\soc/cpu/cpuregs/regs[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5381_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0279_ ),
    .Q(\soc/cpu/cpuregs/regs[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5382_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0280_ ),
    .Q(\soc/cpu/cpuregs/regs[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5383_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0281_ ),
    .Q(\soc/cpu/cpuregs/regs[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5384_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0282_ ),
    .Q(\soc/cpu/cpuregs/regs[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5385_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0283_ ),
    .Q(\soc/cpu/cpuregs/regs[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5386_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0284_ ),
    .Q(\soc/cpu/cpuregs/regs[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5387_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0285_ ),
    .Q(\soc/cpu/cpuregs/regs[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5388_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0286_ ),
    .Q(\soc/cpu/cpuregs/regs[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5389_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0287_ ),
    .Q(\soc/cpu/cpuregs/regs[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5390_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0288_ ),
    .Q(\soc/cpu/cpuregs/regs[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5391_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0289_ ),
    .Q(\soc/cpu/cpuregs/regs[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5392_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0290_ ),
    .Q(\soc/cpu/cpuregs/regs[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5393_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0291_ ),
    .Q(\soc/cpu/cpuregs/regs[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5394_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0292_ ),
    .Q(\soc/cpu/cpuregs/regs[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5395_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0293_ ),
    .Q(\soc/cpu/cpuregs/regs[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5396_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0294_ ),
    .Q(\soc/cpu/cpuregs/regs[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5397_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0295_ ),
    .Q(\soc/cpu/cpuregs/regs[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5398_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0296_ ),
    .Q(\soc/cpu/cpuregs/regs[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5399_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0297_ ),
    .Q(\soc/cpu/cpuregs/regs[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5400_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0298_ ),
    .Q(\soc/cpu/cpuregs/regs[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5401_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0299_ ),
    .Q(\soc/cpu/cpuregs/regs[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5402_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0300_ ),
    .Q(\soc/cpu/cpuregs/regs[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5403_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0301_ ),
    .Q(\soc/cpu/cpuregs/regs[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5404_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0302_ ),
    .Q(\soc/cpu/cpuregs/regs[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5405_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0303_ ),
    .Q(\soc/cpu/cpuregs/regs[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5406_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0304_ ),
    .Q(\soc/cpu/cpuregs/regs[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5407_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0305_ ),
    .Q(\soc/cpu/cpuregs/regs[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5408_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0306_ ),
    .Q(\soc/cpu/cpuregs/regs[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5409_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0307_ ),
    .Q(\soc/cpu/cpuregs/regs[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5410_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0308_ ),
    .Q(\soc/cpu/cpuregs/regs[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5411_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0309_ ),
    .Q(\soc/cpu/cpuregs/regs[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5412_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0310_ ),
    .Q(\soc/cpu/cpuregs/regs[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5413_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0311_ ),
    .Q(\soc/cpu/cpuregs/regs[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5414_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0312_ ),
    .Q(\soc/cpu/cpuregs/regs[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5415_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0313_ ),
    .Q(\soc/cpu/cpuregs/regs[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5416_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0314_ ),
    .Q(\soc/cpu/cpuregs/regs[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5417_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0315_ ),
    .Q(\soc/cpu/cpuregs/regs[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5418_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0316_ ),
    .Q(\soc/cpu/cpuregs/regs[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5419_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0317_ ),
    .Q(\soc/cpu/cpuregs/regs[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5420_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0318_ ),
    .Q(\soc/cpu/cpuregs/regs[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5421_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0319_ ),
    .Q(\soc/cpu/cpuregs/regs[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5422_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0320_ ),
    .Q(\soc/cpu/cpuregs/regs[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5423_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0321_ ),
    .Q(\soc/cpu/cpuregs/regs[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5424_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0322_ ),
    .Q(\soc/cpu/cpuregs/regs[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5425_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0323_ ),
    .Q(\soc/cpu/cpuregs/regs[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5426_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0324_ ),
    .Q(\soc/cpu/cpuregs/regs[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5427_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0325_ ),
    .Q(\soc/cpu/cpuregs/regs[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5428_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0326_ ),
    .Q(\soc/cpu/cpuregs/regs[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5429_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0327_ ),
    .Q(\soc/cpu/cpuregs/regs[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5430_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0328_ ),
    .Q(\soc/cpu/cpuregs/regs[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5431_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0329_ ),
    .Q(\soc/cpu/cpuregs/regs[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5432_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0330_ ),
    .Q(\soc/cpu/cpuregs/regs[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5433_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0331_ ),
    .Q(\soc/cpu/cpuregs/regs[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5434_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0332_ ),
    .Q(\soc/cpu/cpuregs/regs[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5435_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0333_ ),
    .Q(\soc/cpu/cpuregs/regs[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5436_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0334_ ),
    .Q(\soc/cpu/cpuregs/regs[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5437_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0335_ ),
    .Q(\soc/cpu/cpuregs/regs[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5438_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0336_ ),
    .Q(\soc/cpu/cpuregs/regs[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5439_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0337_ ),
    .Q(\soc/cpu/cpuregs/regs[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5440_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0338_ ),
    .Q(\soc/cpu/cpuregs/regs[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5441_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0339_ ),
    .Q(\soc/cpu/cpuregs/regs[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5442_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0340_ ),
    .Q(\soc/cpu/cpuregs/regs[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5443_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0341_ ),
    .Q(\soc/cpu/cpuregs/regs[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5444_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0342_ ),
    .Q(\soc/cpu/cpuregs/regs[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5445_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0343_ ),
    .Q(\soc/cpu/cpuregs/regs[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5446_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0344_ ),
    .Q(\soc/cpu/cpuregs/regs[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5447_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0345_ ),
    .Q(\soc/cpu/cpuregs/regs[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5448_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0346_ ),
    .Q(\soc/cpu/cpuregs/regs[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5449_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0347_ ),
    .Q(\soc/cpu/cpuregs/regs[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5450_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0348_ ),
    .Q(\soc/cpu/cpuregs/regs[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5451_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0349_ ),
    .Q(\soc/cpu/cpuregs/regs[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5452_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0350_ ),
    .Q(\soc/cpu/cpuregs/regs[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5453_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0351_ ),
    .Q(\soc/cpu/cpuregs/regs[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5454_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0352_ ),
    .Q(\soc/cpu/cpuregs/regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5455_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0353_ ),
    .Q(\soc/cpu/cpuregs/regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5456_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0354_ ),
    .Q(\soc/cpu/cpuregs/regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5457_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0355_ ),
    .Q(\soc/cpu/cpuregs/regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5458_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0356_ ),
    .Q(\soc/cpu/cpuregs/regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5459_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0357_ ),
    .Q(\soc/cpu/cpuregs/regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5460_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0358_ ),
    .Q(\soc/cpu/cpuregs/regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5461_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0359_ ),
    .Q(\soc/cpu/cpuregs/regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5462_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0360_ ),
    .Q(\soc/cpu/cpuregs/regs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5463_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0361_ ),
    .Q(\soc/cpu/cpuregs/regs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5464_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0362_ ),
    .Q(\soc/cpu/cpuregs/regs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5465_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0363_ ),
    .Q(\soc/cpu/cpuregs/regs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5466_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0364_ ),
    .Q(\soc/cpu/cpuregs/regs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5467_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0365_ ),
    .Q(\soc/cpu/cpuregs/regs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5468_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0366_ ),
    .Q(\soc/cpu/cpuregs/regs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5469_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0367_ ),
    .Q(\soc/cpu/cpuregs/regs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5470_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0368_ ),
    .Q(\soc/cpu/cpuregs/regs[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5471_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0369_ ),
    .Q(\soc/cpu/cpuregs/regs[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5472_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0370_ ),
    .Q(\soc/cpu/cpuregs/regs[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5473_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0371_ ),
    .Q(\soc/cpu/cpuregs/regs[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5474_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0372_ ),
    .Q(\soc/cpu/cpuregs/regs[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5475_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0373_ ),
    .Q(\soc/cpu/cpuregs/regs[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5476_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0374_ ),
    .Q(\soc/cpu/cpuregs/regs[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5477_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0375_ ),
    .Q(\soc/cpu/cpuregs/regs[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5478_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0376_ ),
    .Q(\soc/cpu/cpuregs/regs[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5479_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0377_ ),
    .Q(\soc/cpu/cpuregs/regs[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5480_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/cpuregs/_0378_ ),
    .Q(\soc/cpu/cpuregs/regs[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5481_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0379_ ),
    .Q(\soc/cpu/cpuregs/regs[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5482_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0380_ ),
    .Q(\soc/cpu/cpuregs/regs[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5483_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0381_ ),
    .Q(\soc/cpu/cpuregs/regs[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5484_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0382_ ),
    .Q(\soc/cpu/cpuregs/regs[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5485_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0383_ ),
    .Q(\soc/cpu/cpuregs/regs[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5486_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0384_ ),
    .Q(\soc/cpu/cpuregs/regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5487_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0385_ ),
    .Q(\soc/cpu/cpuregs/regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5488_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0386_ ),
    .Q(\soc/cpu/cpuregs/regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5489_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0387_ ),
    .Q(\soc/cpu/cpuregs/regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5490_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0388_ ),
    .Q(\soc/cpu/cpuregs/regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5491_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0389_ ),
    .Q(\soc/cpu/cpuregs/regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5492_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0390_ ),
    .Q(\soc/cpu/cpuregs/regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5493_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0391_ ),
    .Q(\soc/cpu/cpuregs/regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5494_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0392_ ),
    .Q(\soc/cpu/cpuregs/regs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5495_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0393_ ),
    .Q(\soc/cpu/cpuregs/regs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5496_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0394_ ),
    .Q(\soc/cpu/cpuregs/regs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5497_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0395_ ),
    .Q(\soc/cpu/cpuregs/regs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5498_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0396_ ),
    .Q(\soc/cpu/cpuregs/regs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5499_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0397_ ),
    .Q(\soc/cpu/cpuregs/regs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5500_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0398_ ),
    .Q(\soc/cpu/cpuregs/regs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5501_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0399_ ),
    .Q(\soc/cpu/cpuregs/regs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5502_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0400_ ),
    .Q(\soc/cpu/cpuregs/regs[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5503_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0401_ ),
    .Q(\soc/cpu/cpuregs/regs[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5504_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0402_ ),
    .Q(\soc/cpu/cpuregs/regs[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5505_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0403_ ),
    .Q(\soc/cpu/cpuregs/regs[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5506_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0404_ ),
    .Q(\soc/cpu/cpuregs/regs[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5507_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0405_ ),
    .Q(\soc/cpu/cpuregs/regs[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5508_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0406_ ),
    .Q(\soc/cpu/cpuregs/regs[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5509_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0407_ ),
    .Q(\soc/cpu/cpuregs/regs[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5510_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0408_ ),
    .Q(\soc/cpu/cpuregs/regs[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5511_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0409_ ),
    .Q(\soc/cpu/cpuregs/regs[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5512_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0410_ ),
    .Q(\soc/cpu/cpuregs/regs[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5513_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0411_ ),
    .Q(\soc/cpu/cpuregs/regs[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5514_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0412_ ),
    .Q(\soc/cpu/cpuregs/regs[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5515_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0413_ ),
    .Q(\soc/cpu/cpuregs/regs[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5516_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0414_ ),
    .Q(\soc/cpu/cpuregs/regs[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5517_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0415_ ),
    .Q(\soc/cpu/cpuregs/regs[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5518_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0416_ ),
    .Q(\soc/cpu/cpuregs/regs[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5519_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0417_ ),
    .Q(\soc/cpu/cpuregs/regs[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5520_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0418_ ),
    .Q(\soc/cpu/cpuregs/regs[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5521_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0419_ ),
    .Q(\soc/cpu/cpuregs/regs[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5522_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0420_ ),
    .Q(\soc/cpu/cpuregs/regs[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5523_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0421_ ),
    .Q(\soc/cpu/cpuregs/regs[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5524_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0422_ ),
    .Q(\soc/cpu/cpuregs/regs[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5525_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0423_ ),
    .Q(\soc/cpu/cpuregs/regs[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5526_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0424_ ),
    .Q(\soc/cpu/cpuregs/regs[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5527_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0425_ ),
    .Q(\soc/cpu/cpuregs/regs[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5528_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0426_ ),
    .Q(\soc/cpu/cpuregs/regs[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5529_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0427_ ),
    .Q(\soc/cpu/cpuregs/regs[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5530_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0428_ ),
    .Q(\soc/cpu/cpuregs/regs[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5531_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0429_ ),
    .Q(\soc/cpu/cpuregs/regs[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5532_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0430_ ),
    .Q(\soc/cpu/cpuregs/regs[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5533_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0431_ ),
    .Q(\soc/cpu/cpuregs/regs[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5534_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0432_ ),
    .Q(\soc/cpu/cpuregs/regs[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5535_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0433_ ),
    .Q(\soc/cpu/cpuregs/regs[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5536_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0434_ ),
    .Q(\soc/cpu/cpuregs/regs[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5537_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0435_ ),
    .Q(\soc/cpu/cpuregs/regs[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5538_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0436_ ),
    .Q(\soc/cpu/cpuregs/regs[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5539_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0437_ ),
    .Q(\soc/cpu/cpuregs/regs[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5540_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0438_ ),
    .Q(\soc/cpu/cpuregs/regs[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5541_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0439_ ),
    .Q(\soc/cpu/cpuregs/regs[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5542_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0440_ ),
    .Q(\soc/cpu/cpuregs/regs[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5543_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0441_ ),
    .Q(\soc/cpu/cpuregs/regs[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5544_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0442_ ),
    .Q(\soc/cpu/cpuregs/regs[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5545_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0443_ ),
    .Q(\soc/cpu/cpuregs/regs[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5546_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0444_ ),
    .Q(\soc/cpu/cpuregs/regs[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5547_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0445_ ),
    .Q(\soc/cpu/cpuregs/regs[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5548_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0446_ ),
    .Q(\soc/cpu/cpuregs/regs[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5549_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0447_ ),
    .Q(\soc/cpu/cpuregs/regs[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5550_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0448_ ),
    .Q(\soc/cpu/cpuregs/regs[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5551_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0449_ ),
    .Q(\soc/cpu/cpuregs/regs[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5552_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0450_ ),
    .Q(\soc/cpu/cpuregs/regs[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5553_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0451_ ),
    .Q(\soc/cpu/cpuregs/regs[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5554_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0452_ ),
    .Q(\soc/cpu/cpuregs/regs[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5555_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0453_ ),
    .Q(\soc/cpu/cpuregs/regs[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5556_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0454_ ),
    .Q(\soc/cpu/cpuregs/regs[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5557_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0455_ ),
    .Q(\soc/cpu/cpuregs/regs[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5558_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0456_ ),
    .Q(\soc/cpu/cpuregs/regs[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5559_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0457_ ),
    .Q(\soc/cpu/cpuregs/regs[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5560_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0458_ ),
    .Q(\soc/cpu/cpuregs/regs[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5561_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0459_ ),
    .Q(\soc/cpu/cpuregs/regs[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5562_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0460_ ),
    .Q(\soc/cpu/cpuregs/regs[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5563_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0461_ ),
    .Q(\soc/cpu/cpuregs/regs[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5564_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0462_ ),
    .Q(\soc/cpu/cpuregs/regs[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5565_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0463_ ),
    .Q(\soc/cpu/cpuregs/regs[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5566_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0464_ ),
    .Q(\soc/cpu/cpuregs/regs[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5567_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0465_ ),
    .Q(\soc/cpu/cpuregs/regs[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5568_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0466_ ),
    .Q(\soc/cpu/cpuregs/regs[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5569_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0467_ ),
    .Q(\soc/cpu/cpuregs/regs[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5570_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0468_ ),
    .Q(\soc/cpu/cpuregs/regs[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5571_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0469_ ),
    .Q(\soc/cpu/cpuregs/regs[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5572_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0470_ ),
    .Q(\soc/cpu/cpuregs/regs[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5573_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0471_ ),
    .Q(\soc/cpu/cpuregs/regs[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5574_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0472_ ),
    .Q(\soc/cpu/cpuregs/regs[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5575_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0473_ ),
    .Q(\soc/cpu/cpuregs/regs[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5576_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0474_ ),
    .Q(\soc/cpu/cpuregs/regs[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5577_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0475_ ),
    .Q(\soc/cpu/cpuregs/regs[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5578_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0476_ ),
    .Q(\soc/cpu/cpuregs/regs[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5579_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0477_ ),
    .Q(\soc/cpu/cpuregs/regs[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5580_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0478_ ),
    .Q(\soc/cpu/cpuregs/regs[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5581_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0479_ ),
    .Q(\soc/cpu/cpuregs/regs[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5582_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0480_ ),
    .Q(\soc/cpu/cpuregs/regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5583_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0481_ ),
    .Q(\soc/cpu/cpuregs/regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5584_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0482_ ),
    .Q(\soc/cpu/cpuregs/regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5585_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0483_ ),
    .Q(\soc/cpu/cpuregs/regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5586_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0484_ ),
    .Q(\soc/cpu/cpuregs/regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5587_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0485_ ),
    .Q(\soc/cpu/cpuregs/regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5588_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0486_ ),
    .Q(\soc/cpu/cpuregs/regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5589_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0487_ ),
    .Q(\soc/cpu/cpuregs/regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5590_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0488_ ),
    .Q(\soc/cpu/cpuregs/regs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5591_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0489_ ),
    .Q(\soc/cpu/cpuregs/regs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5592_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0490_ ),
    .Q(\soc/cpu/cpuregs/regs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5593_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0491_ ),
    .Q(\soc/cpu/cpuregs/regs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5594_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0492_ ),
    .Q(\soc/cpu/cpuregs/regs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5595_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0493_ ),
    .Q(\soc/cpu/cpuregs/regs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5596_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0494_ ),
    .Q(\soc/cpu/cpuregs/regs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5597_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0495_ ),
    .Q(\soc/cpu/cpuregs/regs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5598_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0496_ ),
    .Q(\soc/cpu/cpuregs/regs[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5599_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0497_ ),
    .Q(\soc/cpu/cpuregs/regs[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5600_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0498_ ),
    .Q(\soc/cpu/cpuregs/regs[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5601_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0499_ ),
    .Q(\soc/cpu/cpuregs/regs[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5602_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0500_ ),
    .Q(\soc/cpu/cpuregs/regs[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5603_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0501_ ),
    .Q(\soc/cpu/cpuregs/regs[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5604_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0502_ ),
    .Q(\soc/cpu/cpuregs/regs[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5605_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0503_ ),
    .Q(\soc/cpu/cpuregs/regs[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5606_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0504_ ),
    .Q(\soc/cpu/cpuregs/regs[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5607_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0505_ ),
    .Q(\soc/cpu/cpuregs/regs[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5608_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0506_ ),
    .Q(\soc/cpu/cpuregs/regs[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5609_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0507_ ),
    .Q(\soc/cpu/cpuregs/regs[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5610_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0508_ ),
    .Q(\soc/cpu/cpuregs/regs[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5611_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0509_ ),
    .Q(\soc/cpu/cpuregs/regs[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5612_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0510_ ),
    .Q(\soc/cpu/cpuregs/regs[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5613_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0511_ ),
    .Q(\soc/cpu/cpuregs/regs[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5614_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0512_ ),
    .Q(\soc/cpu/cpuregs/regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5615_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0513_ ),
    .Q(\soc/cpu/cpuregs/regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5616_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0514_ ),
    .Q(\soc/cpu/cpuregs/regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5617_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0515_ ),
    .Q(\soc/cpu/cpuregs/regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5618_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0516_ ),
    .Q(\soc/cpu/cpuregs/regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5619_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0517_ ),
    .Q(\soc/cpu/cpuregs/regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5620_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0518_ ),
    .Q(\soc/cpu/cpuregs/regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5621_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0519_ ),
    .Q(\soc/cpu/cpuregs/regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5622_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0520_ ),
    .Q(\soc/cpu/cpuregs/regs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5623_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0521_ ),
    .Q(\soc/cpu/cpuregs/regs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5624_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0522_ ),
    .Q(\soc/cpu/cpuregs/regs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5625_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0523_ ),
    .Q(\soc/cpu/cpuregs/regs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5626_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0524_ ),
    .Q(\soc/cpu/cpuregs/regs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5627_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0525_ ),
    .Q(\soc/cpu/cpuregs/regs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5628_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0526_ ),
    .Q(\soc/cpu/cpuregs/regs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5629_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0527_ ),
    .Q(\soc/cpu/cpuregs/regs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5630_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0528_ ),
    .Q(\soc/cpu/cpuregs/regs[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5631_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0529_ ),
    .Q(\soc/cpu/cpuregs/regs[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5632_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0530_ ),
    .Q(\soc/cpu/cpuregs/regs[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5633_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0531_ ),
    .Q(\soc/cpu/cpuregs/regs[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5634_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0532_ ),
    .Q(\soc/cpu/cpuregs/regs[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5635_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0533_ ),
    .Q(\soc/cpu/cpuregs/regs[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5636_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0534_ ),
    .Q(\soc/cpu/cpuregs/regs[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5637_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0535_ ),
    .Q(\soc/cpu/cpuregs/regs[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5638_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0536_ ),
    .Q(\soc/cpu/cpuregs/regs[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5639_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0537_ ),
    .Q(\soc/cpu/cpuregs/regs[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5640_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0538_ ),
    .Q(\soc/cpu/cpuregs/regs[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5641_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0539_ ),
    .Q(\soc/cpu/cpuregs/regs[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5642_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0540_ ),
    .Q(\soc/cpu/cpuregs/regs[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5643_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0541_ ),
    .Q(\soc/cpu/cpuregs/regs[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5644_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0542_ ),
    .Q(\soc/cpu/cpuregs/regs[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5645_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0543_ ),
    .Q(\soc/cpu/cpuregs/regs[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5646_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0544_ ),
    .Q(\soc/cpu/cpuregs/regs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5647_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0545_ ),
    .Q(\soc/cpu/cpuregs/regs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5648_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0546_ ),
    .Q(\soc/cpu/cpuregs/regs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5649_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0547_ ),
    .Q(\soc/cpu/cpuregs/regs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5650_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0548_ ),
    .Q(\soc/cpu/cpuregs/regs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5651_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0549_ ),
    .Q(\soc/cpu/cpuregs/regs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5652_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0550_ ),
    .Q(\soc/cpu/cpuregs/regs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5653_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0551_ ),
    .Q(\soc/cpu/cpuregs/regs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5654_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0552_ ),
    .Q(\soc/cpu/cpuregs/regs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5655_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0553_ ),
    .Q(\soc/cpu/cpuregs/regs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5656_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0554_ ),
    .Q(\soc/cpu/cpuregs/regs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5657_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0555_ ),
    .Q(\soc/cpu/cpuregs/regs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5658_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0556_ ),
    .Q(\soc/cpu/cpuregs/regs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5659_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0557_ ),
    .Q(\soc/cpu/cpuregs/regs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5660_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0558_ ),
    .Q(\soc/cpu/cpuregs/regs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5661_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0559_ ),
    .Q(\soc/cpu/cpuregs/regs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5662_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0560_ ),
    .Q(\soc/cpu/cpuregs/regs[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5663_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0561_ ),
    .Q(\soc/cpu/cpuregs/regs[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5664_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0562_ ),
    .Q(\soc/cpu/cpuregs/regs[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5665_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0563_ ),
    .Q(\soc/cpu/cpuregs/regs[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5666_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0564_ ),
    .Q(\soc/cpu/cpuregs/regs[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5667_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0565_ ),
    .Q(\soc/cpu/cpuregs/regs[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5668_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0566_ ),
    .Q(\soc/cpu/cpuregs/regs[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5669_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0567_ ),
    .Q(\soc/cpu/cpuregs/regs[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5670_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0568_ ),
    .Q(\soc/cpu/cpuregs/regs[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5671_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0569_ ),
    .Q(\soc/cpu/cpuregs/regs[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5672_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0570_ ),
    .Q(\soc/cpu/cpuregs/regs[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5673_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0571_ ),
    .Q(\soc/cpu/cpuregs/regs[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5674_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0572_ ),
    .Q(\soc/cpu/cpuregs/regs[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5675_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0573_ ),
    .Q(\soc/cpu/cpuregs/regs[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5676_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0574_ ),
    .Q(\soc/cpu/cpuregs/regs[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5677_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0575_ ),
    .Q(\soc/cpu/cpuregs/regs[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5678_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0576_ ),
    .Q(\soc/cpu/cpuregs/regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5679_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0577_ ),
    .Q(\soc/cpu/cpuregs/regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5680_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0578_ ),
    .Q(\soc/cpu/cpuregs/regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5681_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0579_ ),
    .Q(\soc/cpu/cpuregs/regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5682_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0580_ ),
    .Q(\soc/cpu/cpuregs/regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5683_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0581_ ),
    .Q(\soc/cpu/cpuregs/regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5684_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0582_ ),
    .Q(\soc/cpu/cpuregs/regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5685_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0583_ ),
    .Q(\soc/cpu/cpuregs/regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5686_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0584_ ),
    .Q(\soc/cpu/cpuregs/regs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5687_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0585_ ),
    .Q(\soc/cpu/cpuregs/regs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5688_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0586_ ),
    .Q(\soc/cpu/cpuregs/regs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5689_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0587_ ),
    .Q(\soc/cpu/cpuregs/regs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5690_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0588_ ),
    .Q(\soc/cpu/cpuregs/regs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5691_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0589_ ),
    .Q(\soc/cpu/cpuregs/regs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5692_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0590_ ),
    .Q(\soc/cpu/cpuregs/regs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5693_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0591_ ),
    .Q(\soc/cpu/cpuregs/regs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5694_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0592_ ),
    .Q(\soc/cpu/cpuregs/regs[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5695_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0593_ ),
    .Q(\soc/cpu/cpuregs/regs[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5696_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0594_ ),
    .Q(\soc/cpu/cpuregs/regs[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5697_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0595_ ),
    .Q(\soc/cpu/cpuregs/regs[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5698_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0596_ ),
    .Q(\soc/cpu/cpuregs/regs[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5699_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0597_ ),
    .Q(\soc/cpu/cpuregs/regs[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5700_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0598_ ),
    .Q(\soc/cpu/cpuregs/regs[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5701_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0599_ ),
    .Q(\soc/cpu/cpuregs/regs[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5702_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0600_ ),
    .Q(\soc/cpu/cpuregs/regs[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5703_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0601_ ),
    .Q(\soc/cpu/cpuregs/regs[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5704_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0602_ ),
    .Q(\soc/cpu/cpuregs/regs[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5705_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0603_ ),
    .Q(\soc/cpu/cpuregs/regs[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5706_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0604_ ),
    .Q(\soc/cpu/cpuregs/regs[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5707_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0605_ ),
    .Q(\soc/cpu/cpuregs/regs[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5708_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0606_ ),
    .Q(\soc/cpu/cpuregs/regs[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5709_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0607_ ),
    .Q(\soc/cpu/cpuregs/regs[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5710_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0608_ ),
    .Q(\soc/cpu/cpuregs/regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5711_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0609_ ),
    .Q(\soc/cpu/cpuregs/regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5712_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0610_ ),
    .Q(\soc/cpu/cpuregs/regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5713_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0611_ ),
    .Q(\soc/cpu/cpuregs/regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5714_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0612_ ),
    .Q(\soc/cpu/cpuregs/regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5715_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0613_ ),
    .Q(\soc/cpu/cpuregs/regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5716_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0614_ ),
    .Q(\soc/cpu/cpuregs/regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5717_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0615_ ),
    .Q(\soc/cpu/cpuregs/regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5718_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0616_ ),
    .Q(\soc/cpu/cpuregs/regs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5719_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0617_ ),
    .Q(\soc/cpu/cpuregs/regs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5720_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0618_ ),
    .Q(\soc/cpu/cpuregs/regs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5721_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0619_ ),
    .Q(\soc/cpu/cpuregs/regs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5722_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0620_ ),
    .Q(\soc/cpu/cpuregs/regs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5723_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0621_ ),
    .Q(\soc/cpu/cpuregs/regs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5724_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0622_ ),
    .Q(\soc/cpu/cpuregs/regs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5725_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0623_ ),
    .Q(\soc/cpu/cpuregs/regs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5726_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0624_ ),
    .Q(\soc/cpu/cpuregs/regs[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5727_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0625_ ),
    .Q(\soc/cpu/cpuregs/regs[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5728_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0626_ ),
    .Q(\soc/cpu/cpuregs/regs[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5729_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0627_ ),
    .Q(\soc/cpu/cpuregs/regs[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5730_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0628_ ),
    .Q(\soc/cpu/cpuregs/regs[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5731_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0629_ ),
    .Q(\soc/cpu/cpuregs/regs[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5732_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0630_ ),
    .Q(\soc/cpu/cpuregs/regs[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5733_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0631_ ),
    .Q(\soc/cpu/cpuregs/regs[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5734_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0632_ ),
    .Q(\soc/cpu/cpuregs/regs[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5735_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0633_ ),
    .Q(\soc/cpu/cpuregs/regs[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5736_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0634_ ),
    .Q(\soc/cpu/cpuregs/regs[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5737_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0635_ ),
    .Q(\soc/cpu/cpuregs/regs[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5738_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0636_ ),
    .Q(\soc/cpu/cpuregs/regs[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5739_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0637_ ),
    .Q(\soc/cpu/cpuregs/regs[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5740_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0638_ ),
    .Q(\soc/cpu/cpuregs/regs[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5741_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0639_ ),
    .Q(\soc/cpu/cpuregs/regs[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5742_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0640_ ),
    .Q(\soc/cpu/cpuregs/regs[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5743_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0641_ ),
    .Q(\soc/cpu/cpuregs/regs[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5744_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0642_ ),
    .Q(\soc/cpu/cpuregs/regs[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5745_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0643_ ),
    .Q(\soc/cpu/cpuregs/regs[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5746_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0644_ ),
    .Q(\soc/cpu/cpuregs/regs[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5747_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0645_ ),
    .Q(\soc/cpu/cpuregs/regs[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5748_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0646_ ),
    .Q(\soc/cpu/cpuregs/regs[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5749_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0647_ ),
    .Q(\soc/cpu/cpuregs/regs[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5750_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0648_ ),
    .Q(\soc/cpu/cpuregs/regs[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5751_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0649_ ),
    .Q(\soc/cpu/cpuregs/regs[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5752_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0650_ ),
    .Q(\soc/cpu/cpuregs/regs[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5753_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0651_ ),
    .Q(\soc/cpu/cpuregs/regs[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5754_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0652_ ),
    .Q(\soc/cpu/cpuregs/regs[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5755_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0653_ ),
    .Q(\soc/cpu/cpuregs/regs[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5756_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0654_ ),
    .Q(\soc/cpu/cpuregs/regs[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5757_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0655_ ),
    .Q(\soc/cpu/cpuregs/regs[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5758_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0656_ ),
    .Q(\soc/cpu/cpuregs/regs[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5759_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0657_ ),
    .Q(\soc/cpu/cpuregs/regs[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5760_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0658_ ),
    .Q(\soc/cpu/cpuregs/regs[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5761_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0659_ ),
    .Q(\soc/cpu/cpuregs/regs[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5762_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0660_ ),
    .Q(\soc/cpu/cpuregs/regs[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5763_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0661_ ),
    .Q(\soc/cpu/cpuregs/regs[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5764_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0662_ ),
    .Q(\soc/cpu/cpuregs/regs[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5765_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0663_ ),
    .Q(\soc/cpu/cpuregs/regs[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5766_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0664_ ),
    .Q(\soc/cpu/cpuregs/regs[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5767_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0665_ ),
    .Q(\soc/cpu/cpuregs/regs[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5768_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0666_ ),
    .Q(\soc/cpu/cpuregs/regs[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5769_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0667_ ),
    .Q(\soc/cpu/cpuregs/regs[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5770_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0668_ ),
    .Q(\soc/cpu/cpuregs/regs[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5771_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0669_ ),
    .Q(\soc/cpu/cpuregs/regs[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5772_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0670_ ),
    .Q(\soc/cpu/cpuregs/regs[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5773_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0671_ ),
    .Q(\soc/cpu/cpuregs/regs[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5774_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0672_ ),
    .Q(\soc/cpu/cpuregs/regs[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5775_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0673_ ),
    .Q(\soc/cpu/cpuregs/regs[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5776_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0674_ ),
    .Q(\soc/cpu/cpuregs/regs[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5777_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0675_ ),
    .Q(\soc/cpu/cpuregs/regs[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5778_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0676_ ),
    .Q(\soc/cpu/cpuregs/regs[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5779_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0677_ ),
    .Q(\soc/cpu/cpuregs/regs[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5780_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0678_ ),
    .Q(\soc/cpu/cpuregs/regs[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5781_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0679_ ),
    .Q(\soc/cpu/cpuregs/regs[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5782_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0680_ ),
    .Q(\soc/cpu/cpuregs/regs[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5783_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0681_ ),
    .Q(\soc/cpu/cpuregs/regs[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5784_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0682_ ),
    .Q(\soc/cpu/cpuregs/regs[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5785_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0683_ ),
    .Q(\soc/cpu/cpuregs/regs[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5786_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0684_ ),
    .Q(\soc/cpu/cpuregs/regs[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5787_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0685_ ),
    .Q(\soc/cpu/cpuregs/regs[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5788_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0686_ ),
    .Q(\soc/cpu/cpuregs/regs[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5789_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0687_ ),
    .Q(\soc/cpu/cpuregs/regs[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5790_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0688_ ),
    .Q(\soc/cpu/cpuregs/regs[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5791_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0689_ ),
    .Q(\soc/cpu/cpuregs/regs[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5792_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0690_ ),
    .Q(\soc/cpu/cpuregs/regs[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5793_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0691_ ),
    .Q(\soc/cpu/cpuregs/regs[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5794_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0692_ ),
    .Q(\soc/cpu/cpuregs/regs[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5795_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0693_ ),
    .Q(\soc/cpu/cpuregs/regs[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5796_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0694_ ),
    .Q(\soc/cpu/cpuregs/regs[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5797_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0695_ ),
    .Q(\soc/cpu/cpuregs/regs[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5798_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0696_ ),
    .Q(\soc/cpu/cpuregs/regs[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5799_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0697_ ),
    .Q(\soc/cpu/cpuregs/regs[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5800_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0698_ ),
    .Q(\soc/cpu/cpuregs/regs[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5801_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0699_ ),
    .Q(\soc/cpu/cpuregs/regs[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5802_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0700_ ),
    .Q(\soc/cpu/cpuregs/regs[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5803_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0701_ ),
    .Q(\soc/cpu/cpuregs/regs[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5804_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0702_ ),
    .Q(\soc/cpu/cpuregs/regs[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5805_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0703_ ),
    .Q(\soc/cpu/cpuregs/regs[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5806_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0704_ ),
    .Q(\soc/cpu/cpuregs/regs[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5807_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0705_ ),
    .Q(\soc/cpu/cpuregs/regs[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5808_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0706_ ),
    .Q(\soc/cpu/cpuregs/regs[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5809_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0707_ ),
    .Q(\soc/cpu/cpuregs/regs[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5810_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0708_ ),
    .Q(\soc/cpu/cpuregs/regs[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5811_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0709_ ),
    .Q(\soc/cpu/cpuregs/regs[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5812_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0710_ ),
    .Q(\soc/cpu/cpuregs/regs[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5813_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0711_ ),
    .Q(\soc/cpu/cpuregs/regs[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5814_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0712_ ),
    .Q(\soc/cpu/cpuregs/regs[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5815_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0713_ ),
    .Q(\soc/cpu/cpuregs/regs[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5816_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0714_ ),
    .Q(\soc/cpu/cpuregs/regs[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5817_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0715_ ),
    .Q(\soc/cpu/cpuregs/regs[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5818_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0716_ ),
    .Q(\soc/cpu/cpuregs/regs[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5819_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0717_ ),
    .Q(\soc/cpu/cpuregs/regs[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5820_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0718_ ),
    .Q(\soc/cpu/cpuregs/regs[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5821_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0719_ ),
    .Q(\soc/cpu/cpuregs/regs[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5822_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0720_ ),
    .Q(\soc/cpu/cpuregs/regs[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5823_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0721_ ),
    .Q(\soc/cpu/cpuregs/regs[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5824_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0722_ ),
    .Q(\soc/cpu/cpuregs/regs[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5825_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0723_ ),
    .Q(\soc/cpu/cpuregs/regs[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5826_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0724_ ),
    .Q(\soc/cpu/cpuregs/regs[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5827_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0725_ ),
    .Q(\soc/cpu/cpuregs/regs[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5828_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0726_ ),
    .Q(\soc/cpu/cpuregs/regs[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5829_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0727_ ),
    .Q(\soc/cpu/cpuregs/regs[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5830_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0728_ ),
    .Q(\soc/cpu/cpuregs/regs[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5831_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0729_ ),
    .Q(\soc/cpu/cpuregs/regs[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5832_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/cpuregs/_0730_ ),
    .Q(\soc/cpu/cpuregs/regs[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5833_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0731_ ),
    .Q(\soc/cpu/cpuregs/regs[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5834_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0732_ ),
    .Q(\soc/cpu/cpuregs/regs[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5835_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0733_ ),
    .Q(\soc/cpu/cpuregs/regs[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5836_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0734_ ),
    .Q(\soc/cpu/cpuregs/regs[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5837_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0735_ ),
    .Q(\soc/cpu/cpuregs/regs[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5838_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0736_ ),
    .Q(\soc/cpu/cpuregs/regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5839_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0737_ ),
    .Q(\soc/cpu/cpuregs/regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5840_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0738_ ),
    .Q(\soc/cpu/cpuregs/regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5841_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0739_ ),
    .Q(\soc/cpu/cpuregs/regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5842_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0740_ ),
    .Q(\soc/cpu/cpuregs/regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5843_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0741_ ),
    .Q(\soc/cpu/cpuregs/regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5844_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0742_ ),
    .Q(\soc/cpu/cpuregs/regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5845_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0743_ ),
    .Q(\soc/cpu/cpuregs/regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5846_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0744_ ),
    .Q(\soc/cpu/cpuregs/regs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5847_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0745_ ),
    .Q(\soc/cpu/cpuregs/regs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5848_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0746_ ),
    .Q(\soc/cpu/cpuregs/regs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5849_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0747_ ),
    .Q(\soc/cpu/cpuregs/regs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5850_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0748_ ),
    .Q(\soc/cpu/cpuregs/regs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5851_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0749_ ),
    .Q(\soc/cpu/cpuregs/regs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5852_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0750_ ),
    .Q(\soc/cpu/cpuregs/regs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5853_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0751_ ),
    .Q(\soc/cpu/cpuregs/regs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5854_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0752_ ),
    .Q(\soc/cpu/cpuregs/regs[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5855_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0753_ ),
    .Q(\soc/cpu/cpuregs/regs[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5856_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0754_ ),
    .Q(\soc/cpu/cpuregs/regs[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5857_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0755_ ),
    .Q(\soc/cpu/cpuregs/regs[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5858_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0756_ ),
    .Q(\soc/cpu/cpuregs/regs[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5859_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0757_ ),
    .Q(\soc/cpu/cpuregs/regs[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5860_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0758_ ),
    .Q(\soc/cpu/cpuregs/regs[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5861_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0759_ ),
    .Q(\soc/cpu/cpuregs/regs[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5862_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0760_ ),
    .Q(\soc/cpu/cpuregs/regs[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5863_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0761_ ),
    .Q(\soc/cpu/cpuregs/regs[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5864_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0762_ ),
    .Q(\soc/cpu/cpuregs/regs[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5865_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0763_ ),
    .Q(\soc/cpu/cpuregs/regs[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5866_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0764_ ),
    .Q(\soc/cpu/cpuregs/regs[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5867_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0765_ ),
    .Q(\soc/cpu/cpuregs/regs[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5868_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0766_ ),
    .Q(\soc/cpu/cpuregs/regs[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5869_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0767_ ),
    .Q(\soc/cpu/cpuregs/regs[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5870_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0768_ ),
    .Q(\soc/cpu/cpuregs/regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5871_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0769_ ),
    .Q(\soc/cpu/cpuregs/regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5872_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0770_ ),
    .Q(\soc/cpu/cpuregs/regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5873_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0771_ ),
    .Q(\soc/cpu/cpuregs/regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5874_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0772_ ),
    .Q(\soc/cpu/cpuregs/regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5875_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0773_ ),
    .Q(\soc/cpu/cpuregs/regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5876_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0774_ ),
    .Q(\soc/cpu/cpuregs/regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5877_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0775_ ),
    .Q(\soc/cpu/cpuregs/regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5878_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0776_ ),
    .Q(\soc/cpu/cpuregs/regs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5879_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0777_ ),
    .Q(\soc/cpu/cpuregs/regs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5880_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0778_ ),
    .Q(\soc/cpu/cpuregs/regs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5881_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0779_ ),
    .Q(\soc/cpu/cpuregs/regs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5882_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0780_ ),
    .Q(\soc/cpu/cpuregs/regs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5883_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0781_ ),
    .Q(\soc/cpu/cpuregs/regs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5884_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0782_ ),
    .Q(\soc/cpu/cpuregs/regs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5885_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0783_ ),
    .Q(\soc/cpu/cpuregs/regs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5886_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0784_ ),
    .Q(\soc/cpu/cpuregs/regs[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5887_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0785_ ),
    .Q(\soc/cpu/cpuregs/regs[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5888_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0786_ ),
    .Q(\soc/cpu/cpuregs/regs[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5889_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0787_ ),
    .Q(\soc/cpu/cpuregs/regs[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5890_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0788_ ),
    .Q(\soc/cpu/cpuregs/regs[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5891_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0789_ ),
    .Q(\soc/cpu/cpuregs/regs[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5892_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0790_ ),
    .Q(\soc/cpu/cpuregs/regs[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5893_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0791_ ),
    .Q(\soc/cpu/cpuregs/regs[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5894_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0792_ ),
    .Q(\soc/cpu/cpuregs/regs[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5895_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0793_ ),
    .Q(\soc/cpu/cpuregs/regs[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5896_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0794_ ),
    .Q(\soc/cpu/cpuregs/regs[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5897_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0795_ ),
    .Q(\soc/cpu/cpuregs/regs[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5898_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0796_ ),
    .Q(\soc/cpu/cpuregs/regs[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5899_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0797_ ),
    .Q(\soc/cpu/cpuregs/regs[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5900_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0798_ ),
    .Q(\soc/cpu/cpuregs/regs[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5901_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0799_ ),
    .Q(\soc/cpu/cpuregs/regs[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5902_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0800_ ),
    .Q(\soc/cpu/cpuregs/regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5903_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0801_ ),
    .Q(\soc/cpu/cpuregs/regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5904_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0802_ ),
    .Q(\soc/cpu/cpuregs/regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5905_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0803_ ),
    .Q(\soc/cpu/cpuregs/regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5906_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0804_ ),
    .Q(\soc/cpu/cpuregs/regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5907_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0805_ ),
    .Q(\soc/cpu/cpuregs/regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5908_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0806_ ),
    .Q(\soc/cpu/cpuregs/regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5909_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0807_ ),
    .Q(\soc/cpu/cpuregs/regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5910_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0808_ ),
    .Q(\soc/cpu/cpuregs/regs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5911_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0809_ ),
    .Q(\soc/cpu/cpuregs/regs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5912_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0810_ ),
    .Q(\soc/cpu/cpuregs/regs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5913_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0811_ ),
    .Q(\soc/cpu/cpuregs/regs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5914_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0812_ ),
    .Q(\soc/cpu/cpuregs/regs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5915_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0813_ ),
    .Q(\soc/cpu/cpuregs/regs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5916_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0814_ ),
    .Q(\soc/cpu/cpuregs/regs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5917_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0815_ ),
    .Q(\soc/cpu/cpuregs/regs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5918_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0816_ ),
    .Q(\soc/cpu/cpuregs/regs[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5919_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0817_ ),
    .Q(\soc/cpu/cpuregs/regs[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5920_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0818_ ),
    .Q(\soc/cpu/cpuregs/regs[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5921_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0819_ ),
    .Q(\soc/cpu/cpuregs/regs[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5922_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0820_ ),
    .Q(\soc/cpu/cpuregs/regs[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5923_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0821_ ),
    .Q(\soc/cpu/cpuregs/regs[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5924_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0822_ ),
    .Q(\soc/cpu/cpuregs/regs[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5925_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0823_ ),
    .Q(\soc/cpu/cpuregs/regs[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5926_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0824_ ),
    .Q(\soc/cpu/cpuregs/regs[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5927_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0825_ ),
    .Q(\soc/cpu/cpuregs/regs[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5928_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0826_ ),
    .Q(\soc/cpu/cpuregs/regs[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5929_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0827_ ),
    .Q(\soc/cpu/cpuregs/regs[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5930_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0828_ ),
    .Q(\soc/cpu/cpuregs/regs[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5931_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0829_ ),
    .Q(\soc/cpu/cpuregs/regs[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5932_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0830_ ),
    .Q(\soc/cpu/cpuregs/regs[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5933_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0831_ ),
    .Q(\soc/cpu/cpuregs/regs[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5934_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0832_ ),
    .Q(\soc/cpu/cpuregs/regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5935_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0833_ ),
    .Q(\soc/cpu/cpuregs/regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5936_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0834_ ),
    .Q(\soc/cpu/cpuregs/regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5937_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0835_ ),
    .Q(\soc/cpu/cpuregs/regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5938_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0836_ ),
    .Q(\soc/cpu/cpuregs/regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5939_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0837_ ),
    .Q(\soc/cpu/cpuregs/regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5940_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0838_ ),
    .Q(\soc/cpu/cpuregs/regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5941_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0839_ ),
    .Q(\soc/cpu/cpuregs/regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5942_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0840_ ),
    .Q(\soc/cpu/cpuregs/regs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5943_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0841_ ),
    .Q(\soc/cpu/cpuregs/regs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5944_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0842_ ),
    .Q(\soc/cpu/cpuregs/regs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5945_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0843_ ),
    .Q(\soc/cpu/cpuregs/regs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5946_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0844_ ),
    .Q(\soc/cpu/cpuregs/regs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5947_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0845_ ),
    .Q(\soc/cpu/cpuregs/regs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5948_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0846_ ),
    .Q(\soc/cpu/cpuregs/regs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5949_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0847_ ),
    .Q(\soc/cpu/cpuregs/regs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5950_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0848_ ),
    .Q(\soc/cpu/cpuregs/regs[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5951_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0849_ ),
    .Q(\soc/cpu/cpuregs/regs[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5952_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0850_ ),
    .Q(\soc/cpu/cpuregs/regs[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5953_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0851_ ),
    .Q(\soc/cpu/cpuregs/regs[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5954_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0852_ ),
    .Q(\soc/cpu/cpuregs/regs[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5955_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0853_ ),
    .Q(\soc/cpu/cpuregs/regs[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5956_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0854_ ),
    .Q(\soc/cpu/cpuregs/regs[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5957_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0855_ ),
    .Q(\soc/cpu/cpuregs/regs[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5958_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0856_ ),
    .Q(\soc/cpu/cpuregs/regs[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5959_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0857_ ),
    .Q(\soc/cpu/cpuregs/regs[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5960_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0858_ ),
    .Q(\soc/cpu/cpuregs/regs[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5961_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0859_ ),
    .Q(\soc/cpu/cpuregs/regs[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5962_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0860_ ),
    .Q(\soc/cpu/cpuregs/regs[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5963_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0861_ ),
    .Q(\soc/cpu/cpuregs/regs[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5964_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0862_ ),
    .Q(\soc/cpu/cpuregs/regs[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5965_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0863_ ),
    .Q(\soc/cpu/cpuregs/regs[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5966_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0864_ ),
    .Q(\soc/cpu/cpuregs/regs[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5967_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0865_ ),
    .Q(\soc/cpu/cpuregs/regs[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5968_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0866_ ),
    .Q(\soc/cpu/cpuregs/regs[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5969_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0867_ ),
    .Q(\soc/cpu/cpuregs/regs[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5970_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0868_ ),
    .Q(\soc/cpu/cpuregs/regs[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5971_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0869_ ),
    .Q(\soc/cpu/cpuregs/regs[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5972_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0870_ ),
    .Q(\soc/cpu/cpuregs/regs[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5973_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0871_ ),
    .Q(\soc/cpu/cpuregs/regs[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5974_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0872_ ),
    .Q(\soc/cpu/cpuregs/regs[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5975_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0873_ ),
    .Q(\soc/cpu/cpuregs/regs[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5976_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0874_ ),
    .Q(\soc/cpu/cpuregs/regs[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5977_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0875_ ),
    .Q(\soc/cpu/cpuregs/regs[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5978_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0876_ ),
    .Q(\soc/cpu/cpuregs/regs[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5979_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0877_ ),
    .Q(\soc/cpu/cpuregs/regs[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5980_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0878_ ),
    .Q(\soc/cpu/cpuregs/regs[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5981_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0879_ ),
    .Q(\soc/cpu/cpuregs/regs[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5982_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0880_ ),
    .Q(\soc/cpu/cpuregs/regs[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5983_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0881_ ),
    .Q(\soc/cpu/cpuregs/regs[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5984_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0882_ ),
    .Q(\soc/cpu/cpuregs/regs[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5985_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0883_ ),
    .Q(\soc/cpu/cpuregs/regs[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5986_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0884_ ),
    .Q(\soc/cpu/cpuregs/regs[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5987_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0885_ ),
    .Q(\soc/cpu/cpuregs/regs[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5988_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0886_ ),
    .Q(\soc/cpu/cpuregs/regs[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5989_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0887_ ),
    .Q(\soc/cpu/cpuregs/regs[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5990_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0888_ ),
    .Q(\soc/cpu/cpuregs/regs[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5991_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0889_ ),
    .Q(\soc/cpu/cpuregs/regs[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5992_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0890_ ),
    .Q(\soc/cpu/cpuregs/regs[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5993_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0891_ ),
    .Q(\soc/cpu/cpuregs/regs[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5994_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_0892_ ),
    .Q(\soc/cpu/cpuregs/regs[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5995_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0893_ ),
    .Q(\soc/cpu/cpuregs/regs[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5996_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0894_ ),
    .Q(\soc/cpu/cpuregs/regs[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5997_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0895_ ),
    .Q(\soc/cpu/cpuregs/regs[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5998_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0896_ ),
    .Q(\soc/cpu/cpuregs/regs[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_5999_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0897_ ),
    .Q(\soc/cpu/cpuregs/regs[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6000_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0898_ ),
    .Q(\soc/cpu/cpuregs/regs[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6001_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0899_ ),
    .Q(\soc/cpu/cpuregs/regs[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6002_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0900_ ),
    .Q(\soc/cpu/cpuregs/regs[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6003_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0901_ ),
    .Q(\soc/cpu/cpuregs/regs[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6004_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0902_ ),
    .Q(\soc/cpu/cpuregs/regs[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6005_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0903_ ),
    .Q(\soc/cpu/cpuregs/regs[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6006_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0904_ ),
    .Q(\soc/cpu/cpuregs/regs[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6007_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0905_ ),
    .Q(\soc/cpu/cpuregs/regs[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6008_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0906_ ),
    .Q(\soc/cpu/cpuregs/regs[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6009_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0907_ ),
    .Q(\soc/cpu/cpuregs/regs[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6010_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0908_ ),
    .Q(\soc/cpu/cpuregs/regs[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6011_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0909_ ),
    .Q(\soc/cpu/cpuregs/regs[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6012_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0910_ ),
    .Q(\soc/cpu/cpuregs/regs[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6013_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0911_ ),
    .Q(\soc/cpu/cpuregs/regs[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6014_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0912_ ),
    .Q(\soc/cpu/cpuregs/regs[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6015_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0913_ ),
    .Q(\soc/cpu/cpuregs/regs[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6016_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0914_ ),
    .Q(\soc/cpu/cpuregs/regs[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6017_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0915_ ),
    .Q(\soc/cpu/cpuregs/regs[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6018_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0916_ ),
    .Q(\soc/cpu/cpuregs/regs[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6019_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0917_ ),
    .Q(\soc/cpu/cpuregs/regs[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6020_  (.CLK(clknet_leaf_37_clk),
    .D(\soc/cpu/cpuregs/_0918_ ),
    .Q(\soc/cpu/cpuregs/regs[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6021_  (.CLK(clknet_leaf_35_clk),
    .D(\soc/cpu/cpuregs/_0919_ ),
    .Q(\soc/cpu/cpuregs/regs[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6022_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0920_ ),
    .Q(\soc/cpu/cpuregs/regs[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6023_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0921_ ),
    .Q(\soc/cpu/cpuregs/regs[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6024_  (.CLK(clknet_leaf_7_clk),
    .D(\soc/cpu/cpuregs/_0922_ ),
    .Q(\soc/cpu/cpuregs/regs[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6025_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0923_ ),
    .Q(\soc/cpu/cpuregs/regs[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6026_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0924_ ),
    .Q(\soc/cpu/cpuregs/regs[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6027_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0925_ ),
    .Q(\soc/cpu/cpuregs/regs[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6028_  (.CLK(clknet_leaf_50_clk),
    .D(\soc/cpu/cpuregs/_0926_ ),
    .Q(\soc/cpu/cpuregs/regs[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6029_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0927_ ),
    .Q(\soc/cpu/cpuregs/regs[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6030_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0928_ ),
    .Q(\soc/cpu/cpuregs/regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6031_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0929_ ),
    .Q(\soc/cpu/cpuregs/regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6032_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0930_ ),
    .Q(\soc/cpu/cpuregs/regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6033_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0931_ ),
    .Q(\soc/cpu/cpuregs/regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6034_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0932_ ),
    .Q(\soc/cpu/cpuregs/regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6035_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0933_ ),
    .Q(\soc/cpu/cpuregs/regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6036_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0934_ ),
    .Q(\soc/cpu/cpuregs/regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6037_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0935_ ),
    .Q(\soc/cpu/cpuregs/regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6038_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0936_ ),
    .Q(\soc/cpu/cpuregs/regs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6039_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0937_ ),
    .Q(\soc/cpu/cpuregs/regs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6040_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0938_ ),
    .Q(\soc/cpu/cpuregs/regs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6041_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0939_ ),
    .Q(\soc/cpu/cpuregs/regs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6042_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0940_ ),
    .Q(\soc/cpu/cpuregs/regs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6043_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0941_ ),
    .Q(\soc/cpu/cpuregs/regs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6044_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0942_ ),
    .Q(\soc/cpu/cpuregs/regs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6045_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_0943_ ),
    .Q(\soc/cpu/cpuregs/regs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6046_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_0944_ ),
    .Q(\soc/cpu/cpuregs/regs[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6047_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0945_ ),
    .Q(\soc/cpu/cpuregs/regs[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6048_  (.CLK(clknet_leaf_45_clk),
    .D(\soc/cpu/cpuregs/_0946_ ),
    .Q(\soc/cpu/cpuregs/regs[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6049_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0947_ ),
    .Q(\soc/cpu/cpuregs/regs[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6050_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0948_ ),
    .Q(\soc/cpu/cpuregs/regs[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6051_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0949_ ),
    .Q(\soc/cpu/cpuregs/regs[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6052_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0950_ ),
    .Q(\soc/cpu/cpuregs/regs[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6053_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0951_ ),
    .Q(\soc/cpu/cpuregs/regs[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6054_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_0952_ ),
    .Q(\soc/cpu/cpuregs/regs[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6055_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_0953_ ),
    .Q(\soc/cpu/cpuregs/regs[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6056_  (.CLK(clknet_leaf_8_clk),
    .D(\soc/cpu/cpuregs/_0954_ ),
    .Q(\soc/cpu/cpuregs/regs[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6057_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0955_ ),
    .Q(\soc/cpu/cpuregs/regs[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6058_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0956_ ),
    .Q(\soc/cpu/cpuregs/regs[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6059_  (.CLK(clknet_leaf_43_clk),
    .D(\soc/cpu/cpuregs/_0957_ ),
    .Q(\soc/cpu/cpuregs/regs[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6060_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_0958_ ),
    .Q(\soc/cpu/cpuregs/regs[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6061_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0959_ ),
    .Q(\soc/cpu/cpuregs/regs[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6062_  (.CLK(clknet_leaf_29_clk),
    .D(\soc/cpu/cpuregs/_0960_ ),
    .Q(\soc/cpu/cpuregs/regs[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6063_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_0961_ ),
    .Q(\soc/cpu/cpuregs/regs[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6064_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0962_ ),
    .Q(\soc/cpu/cpuregs/regs[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6065_  (.CLK(clknet_leaf_48_clk),
    .D(\soc/cpu/cpuregs/_0963_ ),
    .Q(\soc/cpu/cpuregs/regs[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6066_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0964_ ),
    .Q(\soc/cpu/cpuregs/regs[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6067_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0965_ ),
    .Q(\soc/cpu/cpuregs/regs[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6068_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0966_ ),
    .Q(\soc/cpu/cpuregs/regs[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6069_  (.CLK(clknet_leaf_18_clk),
    .D(\soc/cpu/cpuregs/_0967_ ),
    .Q(\soc/cpu/cpuregs/regs[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6070_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0968_ ),
    .Q(\soc/cpu/cpuregs/regs[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6071_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0969_ ),
    .Q(\soc/cpu/cpuregs/regs[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6072_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0970_ ),
    .Q(\soc/cpu/cpuregs/regs[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6073_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_0971_ ),
    .Q(\soc/cpu/cpuregs/regs[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6074_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0972_ ),
    .Q(\soc/cpu/cpuregs/regs[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6075_  (.CLK(clknet_leaf_17_clk),
    .D(\soc/cpu/cpuregs/_0973_ ),
    .Q(\soc/cpu/cpuregs/regs[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6076_  (.CLK(clknet_leaf_26_clk),
    .D(\soc/cpu/cpuregs/_0974_ ),
    .Q(\soc/cpu/cpuregs/regs[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6077_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0975_ ),
    .Q(\soc/cpu/cpuregs/regs[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6078_  (.CLK(clknet_leaf_12_clk),
    .D(\soc/cpu/cpuregs/_0976_ ),
    .Q(\soc/cpu/cpuregs/regs[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6079_  (.CLK(clknet_leaf_19_clk),
    .D(\soc/cpu/cpuregs/_0977_ ),
    .Q(\soc/cpu/cpuregs/regs[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6080_  (.CLK(clknet_leaf_47_clk),
    .D(\soc/cpu/cpuregs/_0978_ ),
    .Q(\soc/cpu/cpuregs/regs[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6081_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0979_ ),
    .Q(\soc/cpu/cpuregs/regs[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6082_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_0980_ ),
    .Q(\soc/cpu/cpuregs/regs[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6083_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0981_ ),
    .Q(\soc/cpu/cpuregs/regs[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6084_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_0982_ ),
    .Q(\soc/cpu/cpuregs/regs[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6085_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_0983_ ),
    .Q(\soc/cpu/cpuregs/regs[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6086_  (.CLK(clknet_leaf_46_clk),
    .D(\soc/cpu/cpuregs/_0984_ ),
    .Q(\soc/cpu/cpuregs/regs[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6087_  (.CLK(clknet_leaf_24_clk),
    .D(\soc/cpu/cpuregs/_0985_ ),
    .Q(\soc/cpu/cpuregs/regs[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6088_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_0986_ ),
    .Q(\soc/cpu/cpuregs/regs[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6089_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_0987_ ),
    .Q(\soc/cpu/cpuregs/regs[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6090_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_0988_ ),
    .Q(\soc/cpu/cpuregs/regs[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6091_  (.CLK(clknet_leaf_42_clk),
    .D(\soc/cpu/cpuregs/_0989_ ),
    .Q(\soc/cpu/cpuregs/regs[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6092_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0990_ ),
    .Q(\soc/cpu/cpuregs/regs[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6093_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0991_ ),
    .Q(\soc/cpu/cpuregs/regs[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6094_  (.CLK(clknet_leaf_30_clk),
    .D(\soc/cpu/cpuregs/_0992_ ),
    .Q(\soc/cpu/cpuregs/regs[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6095_  (.CLK(clknet_leaf_28_clk),
    .D(\soc/cpu/cpuregs/_0993_ ),
    .Q(\soc/cpu/cpuregs/regs[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6096_  (.CLK(clknet_leaf_49_clk),
    .D(\soc/cpu/cpuregs/_0994_ ),
    .Q(\soc/cpu/cpuregs/regs[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6097_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_0995_ ),
    .Q(\soc/cpu/cpuregs/regs[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6098_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_0996_ ),
    .Q(\soc/cpu/cpuregs/regs[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6099_  (.CLK(clknet_leaf_32_clk),
    .D(\soc/cpu/cpuregs/_0997_ ),
    .Q(\soc/cpu/cpuregs/regs[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6100_  (.CLK(clknet_leaf_16_clk),
    .D(\soc/cpu/cpuregs/_0998_ ),
    .Q(\soc/cpu/cpuregs/regs[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6101_  (.CLK(clknet_leaf_23_clk),
    .D(\soc/cpu/cpuregs/_0999_ ),
    .Q(\soc/cpu/cpuregs/regs[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6102_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_1000_ ),
    .Q(\soc/cpu/cpuregs/regs[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6103_  (.CLK(clknet_leaf_14_clk),
    .D(\soc/cpu/cpuregs/_1001_ ),
    .Q(\soc/cpu/cpuregs/regs[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6104_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_1002_ ),
    .Q(\soc/cpu/cpuregs/regs[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6105_  (.CLK(clknet_leaf_21_clk),
    .D(\soc/cpu/cpuregs/_1003_ ),
    .Q(\soc/cpu/cpuregs/regs[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6106_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_1004_ ),
    .Q(\soc/cpu/cpuregs/regs[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6107_  (.CLK(clknet_leaf_15_clk),
    .D(\soc/cpu/cpuregs/_1005_ ),
    .Q(\soc/cpu/cpuregs/regs[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6108_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_1006_ ),
    .Q(\soc/cpu/cpuregs/regs[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6109_  (.CLK(clknet_leaf_25_clk),
    .D(\soc/cpu/cpuregs/_1007_ ),
    .Q(\soc/cpu/cpuregs/regs[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6110_  (.CLK(clknet_leaf_13_clk),
    .D(\soc/cpu/cpuregs/_1008_ ),
    .Q(\soc/cpu/cpuregs/regs[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6111_  (.CLK(clknet_leaf_20_clk),
    .D(\soc/cpu/cpuregs/_1009_ ),
    .Q(\soc/cpu/cpuregs/regs[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6112_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_1010_ ),
    .Q(\soc/cpu/cpuregs/regs[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6113_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_1011_ ),
    .Q(\soc/cpu/cpuregs/regs[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6114_  (.CLK(clknet_leaf_27_clk),
    .D(\soc/cpu/cpuregs/_1012_ ),
    .Q(\soc/cpu/cpuregs/regs[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6115_  (.CLK(clknet_leaf_52_clk),
    .D(\soc/cpu/cpuregs/_1013_ ),
    .Q(\soc/cpu/cpuregs/regs[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6116_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_1014_ ),
    .Q(\soc/cpu/cpuregs/regs[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6117_  (.CLK(clknet_leaf_33_clk),
    .D(\soc/cpu/cpuregs/_1015_ ),
    .Q(\soc/cpu/cpuregs/regs[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6118_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_1016_ ),
    .Q(\soc/cpu/cpuregs/regs[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6119_  (.CLK(clknet_leaf_22_clk),
    .D(\soc/cpu/cpuregs/_1017_ ),
    .Q(\soc/cpu/cpuregs/regs[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6120_  (.CLK(clknet_leaf_36_clk),
    .D(\soc/cpu/cpuregs/_1018_ ),
    .Q(\soc/cpu/cpuregs/regs[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6121_  (.CLK(clknet_leaf_34_clk),
    .D(\soc/cpu/cpuregs/_1019_ ),
    .Q(\soc/cpu/cpuregs/regs[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6122_  (.CLK(clknet_leaf_38_clk),
    .D(\soc/cpu/cpuregs/_1020_ ),
    .Q(\soc/cpu/cpuregs/regs[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6123_  (.CLK(clknet_leaf_44_clk),
    .D(\soc/cpu/cpuregs/_1021_ ),
    .Q(\soc/cpu/cpuregs/regs[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6124_  (.CLK(clknet_leaf_51_clk),
    .D(\soc/cpu/cpuregs/_1022_ ),
    .Q(\soc/cpu/cpuregs/regs[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/cpu/cpuregs/_6125_  (.CLK(clknet_leaf_31_clk),
    .D(\soc/cpu/cpuregs/_1023_ ),
    .Q(\soc/cpu/cpuregs/regs[16][31] ));
 sram22_256x32m4w8 \soc/memory  (.clk(clknet_leaf_92_clk),
    .we(net495),
    .addr({net525,
    net519,
    net498,
    net509,
    net503,
    net375,
    net382,
    net389}),
    .din({net590,
    net610,
    net168,
    net626,
    net634,
    net646,
    net573,
    net638,
    net587,
    net642,
    net194,
    net618,
    net201,
    net622,
    net630,
    net211,
    net215,
    net582,
    net222,
    net226,
    net230,
    net601,
    net236,
    net243,
    net607,
    net254,
    net593,
    net604,
    net614,
    net269,
    net277,
    net284}),
    .dout({\soc/ram_rdata[31] ,
    \soc/ram_rdata[30] ,
    \soc/ram_rdata[29] ,
    \soc/ram_rdata[28] ,
    \soc/ram_rdata[27] ,
    \soc/ram_rdata[26] ,
    \soc/ram_rdata[25] ,
    \soc/ram_rdata[24] ,
    \soc/ram_rdata[23] ,
    \soc/ram_rdata[22] ,
    \soc/ram_rdata[21] ,
    \soc/ram_rdata[20] ,
    \soc/ram_rdata[19] ,
    \soc/ram_rdata[18] ,
    \soc/ram_rdata[17] ,
    \soc/ram_rdata[16] ,
    \soc/ram_rdata[15] ,
    \soc/ram_rdata[14] ,
    \soc/ram_rdata[13] ,
    \soc/ram_rdata[12] ,
    \soc/ram_rdata[11] ,
    \soc/ram_rdata[10] ,
    \soc/ram_rdata[9] ,
    \soc/ram_rdata[8] ,
    \soc/ram_rdata[7] ,
    \soc/ram_rdata[6] ,
    \soc/ram_rdata[5] ,
    \soc/ram_rdata[4] ,
    \soc/ram_rdata[3] ,
    \soc/ram_rdata[2] ,
    \soc/ram_rdata[1] ,
    \soc/ram_rdata[0] }),
    .wmask({net397,
    net578,
    net564,
    net569}));
 sky130_fd_sc_hd__or3_2 \soc/simpleuart/_0673_  (.A(\soc/simpleuart/send_bitcnt[1] ),
    .B(\soc/simpleuart/send_bitcnt[0] ),
    .C(\soc/simpleuart/send_bitcnt[2] ),
    .X(\soc/simpleuart/_0133_ ));
 sky130_fd_sc_hd__o31a_1 \soc/simpleuart/_0674_  (.A1(\soc/simpleuart/send_bitcnt[3] ),
    .A2(net772),
    .A3(\soc/simpleuart/_0133_ ),
    .B1(\soc/_012_ ),
    .X(\soc/simpleuart_reg_dat_wait ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0675_  (.A(\soc/simpleuart/recv_buf_data[0] ),
    .Y(\soc/simpleuart/_0134_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0677_  (.A(\soc/simpleuart/_0134_ ),
    .B(\soc/simpleuart/recv_buf_valid ),
    .Y(\soc/simpleuart_reg_dat_do[0] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0678_  (.A(\soc/simpleuart/recv_buf_data[1] ),
    .Y(\soc/simpleuart/_0136_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0679_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0136_ ),
    .Y(\soc/simpleuart_reg_dat_do[1] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0680_  (.A(\soc/simpleuart/recv_buf_data[2] ),
    .Y(\soc/simpleuart/_0137_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0681_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0137_ ),
    .Y(\soc/simpleuart_reg_dat_do[2] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0682_  (.A(\soc/simpleuart/recv_buf_data[3] ),
    .Y(\soc/simpleuart/_0138_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0683_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0138_ ),
    .Y(\soc/simpleuart_reg_dat_do[3] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0684_  (.A(\soc/simpleuart/recv_buf_data[4] ),
    .Y(\soc/simpleuart/_0139_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0685_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0139_ ),
    .Y(\soc/simpleuart_reg_dat_do[4] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0686_  (.A(\soc/simpleuart/recv_buf_data[5] ),
    .Y(\soc/simpleuart/_0140_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0687_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0140_ ),
    .Y(\soc/simpleuart_reg_dat_do[5] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0688_  (.A(\soc/simpleuart/recv_buf_data[6] ),
    .Y(\soc/simpleuart/_0141_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0689_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0141_ ),
    .Y(\soc/simpleuart_reg_dat_do[6] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0690_  (.A(\soc/simpleuart/recv_buf_data[7] ),
    .Y(\soc/simpleuart/_0142_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0691_  (.A(\soc/simpleuart/recv_buf_valid ),
    .B(\soc/simpleuart/_0142_ ),
    .Y(\soc/simpleuart_reg_dat_do[7] ));
 sky130_fd_sc_hd__clkinv_8 \soc/simpleuart/_0692_  (.A(\soc/simpleuart/recv_buf_valid ),
    .Y(\soc/simpleuart_reg_dat_do[31] ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0693_  (.A(\soc/simpleuart_reg_div_do[5] ),
    .Y(\soc/simpleuart/_0143_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_0694_  (.A(\soc/simpleuart/send_divcnt[4] ),
    .SLEEP(\soc/simpleuart_reg_div_do[4] ),
    .X(\soc/simpleuart/_0144_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0695_  (.A(\soc/simpleuart_reg_div_do[2] ),
    .Y(\soc/simpleuart/_0145_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0696_  (.A(\soc/simpleuart_reg_div_do[1] ),
    .Y(\soc/simpleuart/_0146_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_0697_  (.A(\soc/simpleuart/send_divcnt[0] ),
    .SLEEP(\soc/simpleuart_reg_div_do[0] ),
    .X(\soc/simpleuart/_0147_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0698_  (.A(\soc/simpleuart/_0146_ ),
    .B(\soc/simpleuart/send_divcnt[1] ),
    .C(\soc/simpleuart/_0147_ ),
    .X(\soc/simpleuart/_0148_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0699_  (.A1(\soc/simpleuart/_0145_ ),
    .A2(\soc/simpleuart/send_divcnt[2] ),
    .B1(\soc/simpleuart/_0148_ ),
    .Y(\soc/simpleuart/_0149_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0700_  (.A(\soc/simpleuart_reg_div_do[3] ),
    .Y(\soc/simpleuart/_0150_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/simpleuart/_0701_  (.A1(\soc/simpleuart/_0150_ ),
    .A2(\soc/simpleuart/send_divcnt[3] ),
    .B1(\soc/simpleuart/send_divcnt[2] ),
    .B2(\soc/simpleuart/_0145_ ),
    .Y(\soc/simpleuart/_0151_ ));
 sky130_fd_sc_hd__clkinv_2 \soc/simpleuart/_0702_  (.A(\soc/simpleuart_reg_div_do[4] ),
    .Y(\soc/simpleuart/_0152_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_0703_  (.A1(\soc/simpleuart/_0152_ ),
    .A2(\soc/simpleuart/send_divcnt[4] ),
    .B1(\soc/simpleuart/send_divcnt[3] ),
    .B2(\soc/simpleuart/_0150_ ),
    .Y(\soc/simpleuart/_0153_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0704_  (.A1(\soc/simpleuart/_0149_ ),
    .A2(\soc/simpleuart/_0151_ ),
    .B1(\soc/simpleuart/_0153_ ),
    .Y(\soc/simpleuart/_0154_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_0705_  (.A1(\soc/simpleuart/_0143_ ),
    .A2(\soc/simpleuart/send_divcnt[5] ),
    .B1(\soc/simpleuart/_0144_ ),
    .B2(\soc/simpleuart/_0154_ ),
    .Y(\soc/simpleuart/_0155_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0706_  (.A(\soc/simpleuart_reg_div_do[6] ),
    .Y(\soc/simpleuart/_0156_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0707_  (.A(\soc/simpleuart/_0156_ ),
    .B(\soc/simpleuart/send_divcnt[6] ),
    .Y(\soc/simpleuart/_0157_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0708_  (.A(\soc/simpleuart/_0143_ ),
    .B(\soc/simpleuart/send_divcnt[5] ),
    .Y(\soc/simpleuart/_0158_ ));
 sky130_fd_sc_hd__inv_2 \soc/simpleuart/_0709_  (.A(\soc/simpleuart_reg_div_do[7] ),
    .Y(\soc/simpleuart/_0159_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_0710_  (.A1(\soc/simpleuart/_0159_ ),
    .A2(\soc/simpleuart/send_divcnt[7] ),
    .B1(\soc/simpleuart/send_divcnt[6] ),
    .B2(\soc/simpleuart/_0156_ ),
    .Y(\soc/simpleuart/_0160_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/simpleuart/_0711_  (.A1(\soc/simpleuart/_0155_ ),
    .A2(\soc/simpleuart/_0157_ ),
    .A3(\soc/simpleuart/_0158_ ),
    .B1(\soc/simpleuart/_0160_ ),
    .Y(\soc/simpleuart/_0161_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0712_  (.A_N(\soc/simpleuart/send_divcnt[8] ),
    .B(\soc/simpleuart_reg_div_do[8] ),
    .Y(\soc/simpleuart/_0162_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0713_  (.A(\soc/simpleuart_reg_div_do[9] ),
    .B(\soc/simpleuart/send_divcnt[9] ),
    .Y(\soc/simpleuart/_0163_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0714_  (.A(\soc/simpleuart/_0159_ ),
    .B(\soc/simpleuart/send_divcnt[7] ),
    .Y(\soc/simpleuart/_0164_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0715_  (.A(\soc/simpleuart_reg_div_do[8] ),
    .Y(\soc/simpleuart/_0165_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0716_  (.A(\soc/simpleuart_reg_div_do[10] ),
    .B(\soc/simpleuart/send_divcnt[10] ),
    .X(\soc/simpleuart/_0166_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0717_  (.A(\soc/simpleuart_reg_div_do[11] ),
    .B(\soc/simpleuart/send_divcnt[11] ),
    .X(\soc/simpleuart/_0167_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/simpleuart/_0718_  (.A1(\soc/simpleuart/_0165_ ),
    .A2(\soc/simpleuart/send_divcnt[8] ),
    .B1(\soc/simpleuart/_0166_ ),
    .C1(\soc/simpleuart/_0167_ ),
    .Y(\soc/simpleuart/_0168_ ));
 sky130_fd_sc_hd__nand4_1 \soc/simpleuart/_0719_  (.A(\soc/simpleuart/_0162_ ),
    .B(\soc/simpleuart/_0163_ ),
    .C(\soc/simpleuart/_0164_ ),
    .D(\soc/simpleuart/_0168_ ),
    .Y(\soc/simpleuart/_0169_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0720_  (.A(\soc/simpleuart_reg_div_do[9] ),
    .Y(\soc/simpleuart/_0170_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0721_  (.A(\soc/simpleuart/_0170_ ),
    .B(\soc/simpleuart/send_divcnt[9] ),
    .C(\soc/simpleuart/_0162_ ),
    .X(\soc/simpleuart/_0171_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0722_  (.A(\soc/simpleuart_reg_div_do[11] ),
    .Y(\soc/simpleuart/_0172_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0723_  (.A_N(\soc/simpleuart/send_divcnt[10] ),
    .B(\soc/simpleuart_reg_div_do[10] ),
    .Y(\soc/simpleuart/_0173_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0724_  (.A(\soc/simpleuart/_0172_ ),
    .B(\soc/simpleuart/send_divcnt[11] ),
    .C(\soc/simpleuart/_0173_ ),
    .X(\soc/simpleuart/_0174_ ));
 sky130_fd_sc_hd__o31a_1 \soc/simpleuart/_0725_  (.A1(\soc/simpleuart/_0166_ ),
    .A2(\soc/simpleuart/_0167_ ),
    .A3(\soc/simpleuart/_0171_ ),
    .B1(\soc/simpleuart/_0174_ ),
    .X(\soc/simpleuart/_0175_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/simpleuart/_0726_  (.A1(\soc/simpleuart/_0161_ ),
    .A2(\soc/simpleuart/_0169_ ),
    .B1(\soc/simpleuart/_0175_ ),
    .Y(\soc/simpleuart/_0176_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0727_  (.A(\soc/simpleuart_reg_div_do[12] ),
    .Y(\soc/simpleuart/_0177_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0728_  (.A(\soc/simpleuart_reg_div_do[13] ),
    .Y(\soc/simpleuart/_0178_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0729_  (.A(\soc/simpleuart/_0178_ ),
    .B(\soc/simpleuart/send_divcnt[13] ),
    .Y(\soc/simpleuart/_0179_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0730_  (.A1(\soc/simpleuart/_0177_ ),
    .A2(\soc/simpleuart/send_divcnt[12] ),
    .B1(\soc/simpleuart/_0179_ ),
    .Y(\soc/simpleuart/_0180_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0731_  (.A(\soc/simpleuart_reg_div_do[14] ),
    .B(\soc/simpleuart/send_divcnt[14] ),
    .X(\soc/simpleuart/_0181_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0732_  (.A(\soc/simpleuart_reg_div_do[15] ),
    .B(\soc/simpleuart/send_divcnt[15] ),
    .X(\soc/simpleuart/_0182_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0733_  (.A(\soc/simpleuart/_0177_ ),
    .B(\soc/simpleuart/send_divcnt[12] ),
    .Y(\soc/simpleuart/_0183_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0734_  (.A(\soc/simpleuart/_0178_ ),
    .B(\soc/simpleuart/send_divcnt[13] ),
    .Y(\soc/simpleuart/_0184_ ));
 sky130_fd_sc_hd__nor4b_1 \soc/simpleuart/_0735_  (.A(\soc/simpleuart/_0181_ ),
    .B(\soc/simpleuart/_0182_ ),
    .C(\soc/simpleuart/_0183_ ),
    .D_N(\soc/simpleuart/_0184_ ),
    .Y(\soc/simpleuart/_0185_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0736_  (.A1(\soc/simpleuart/_0183_ ),
    .A2(\soc/simpleuart/_0184_ ),
    .B1(\soc/simpleuart/_0179_ ),
    .Y(\soc/simpleuart/_0186_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0737_  (.A(\soc/simpleuart_reg_div_do[15] ),
    .Y(\soc/simpleuart/_0187_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0738_  (.A_N(\soc/simpleuart/send_divcnt[14] ),
    .B(\soc/simpleuart_reg_div_do[14] ),
    .Y(\soc/simpleuart/_0188_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0739_  (.A(\soc/simpleuart/_0187_ ),
    .B(\soc/simpleuart/send_divcnt[15] ),
    .C(\soc/simpleuart/_0188_ ),
    .X(\soc/simpleuart/_0189_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/simpleuart/_0740_  (.A1(\soc/simpleuart/_0181_ ),
    .A2(\soc/simpleuart/_0182_ ),
    .A3(\soc/simpleuart/_0186_ ),
    .B1(\soc/simpleuart/_0189_ ),
    .Y(\soc/simpleuart/_0190_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/simpleuart/_0741_  (.A1(\soc/simpleuart/_0176_ ),
    .A2(\soc/simpleuart/_0180_ ),
    .A3(\soc/simpleuart/_0185_ ),
    .B1(\soc/simpleuart/_0190_ ),
    .Y(\soc/simpleuart/_0191_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0742_  (.A(\soc/simpleuart_reg_div_do[26] ),
    .Y(\soc/simpleuart/_0192_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0743_  (.A(\soc/simpleuart_reg_div_do[27] ),
    .Y(\soc/simpleuart/_0193_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0744_  (.A_N(\soc/simpleuart/send_divcnt[26] ),
    .B(\soc/simpleuart_reg_div_do[26] ),
    .Y(\soc/simpleuart/_0194_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0745_  (.A1(\soc/simpleuart/_0193_ ),
    .A2(\soc/simpleuart/send_divcnt[27] ),
    .B1(\soc/simpleuart/_0194_ ),
    .Y(\soc/simpleuart/_0195_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_0746_  (.A(\soc/simpleuart/send_divcnt[27] ),
    .SLEEP(\soc/simpleuart_reg_div_do[27] ),
    .X(\soc/simpleuart/_0196_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/simpleuart/_0747_  (.A1(\soc/simpleuart/_0192_ ),
    .A2(\soc/simpleuart/send_divcnt[26] ),
    .B1(\soc/simpleuart/_0195_ ),
    .C1(\soc/simpleuart/_0196_ ),
    .Y(\soc/simpleuart/_0197_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0748_  (.A(\soc/simpleuart/send_divcnt[24] ),
    .Y(\soc/simpleuart/_0198_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0749_  (.A(\soc/simpleuart_reg_div_do[24] ),
    .B(\soc/simpleuart/_0198_ ),
    .Y(\soc/simpleuart/_0199_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0750_  (.A_N(\soc/simpleuart/send_divcnt[25] ),
    .B(\soc/simpleuart_reg_div_do[25] ),
    .Y(\soc/simpleuart/_0200_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0751_  (.A1(\soc/simpleuart_reg_div_do[24] ),
    .A2(\soc/simpleuart/_0198_ ),
    .B1(\soc/simpleuart/_0200_ ),
    .Y(\soc/simpleuart/_0201_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_0752_  (.A(\soc/simpleuart/send_divcnt[25] ),
    .SLEEP(\soc/simpleuart_reg_div_do[25] ),
    .X(\soc/simpleuart/_0202_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0753_  (.A(\soc/simpleuart/_0201_ ),
    .B(\soc/simpleuart/_0202_ ),
    .Y(\soc/simpleuart/_0203_ ));
 sky130_fd_sc_hd__nand3_2 \soc/simpleuart/_0754_  (.A(\soc/simpleuart/_0197_ ),
    .B(\soc/simpleuart/_0199_ ),
    .C(\soc/simpleuart/_0203_ ),
    .Y(\soc/simpleuart/_0204_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0755_  (.A(\soc/simpleuart/send_divcnt[29] ),
    .Y(\soc/simpleuart/_0205_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_0756_  (.A(\soc/simpleuart_reg_div_do[31] ),
    .SLEEP(\soc/simpleuart/send_divcnt[31] ),
    .X(\soc/simpleuart/_0206_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_0757_  (.A(\soc/simpleuart/send_divcnt[31] ),
    .SLEEP(\soc/simpleuart_reg_div_do[31] ),
    .X(\soc/simpleuart/_0207_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0758_  (.A(\soc/simpleuart_reg_div_do[30] ),
    .B(\soc/simpleuart/send_divcnt[30] ),
    .X(\soc/simpleuart/_0208_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0759_  (.A(\soc/simpleuart/_0206_ ),
    .B(\soc/simpleuart/_0207_ ),
    .C(\soc/simpleuart/_0208_ ),
    .Y(\soc/simpleuart/_0209_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_0760_  (.A1(\soc/simpleuart_reg_div_do[29] ),
    .A2(\soc/simpleuart/_0205_ ),
    .B1(\soc/simpleuart/_0209_ ),
    .Y(\soc/simpleuart/_0210_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0761_  (.A(\soc/simpleuart/send_divcnt[28] ),
    .Y(\soc/simpleuart/_0211_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/simpleuart/_0762_  (.A1(\soc/simpleuart_reg_div_do[29] ),
    .A2(\soc/simpleuart/_0205_ ),
    .B1(\soc/simpleuart/_0211_ ),
    .B2(\soc/simpleuart_reg_div_do[28] ),
    .Y(\soc/simpleuart/_0212_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0763_  (.A1(\soc/simpleuart_reg_div_do[28] ),
    .A2(\soc/simpleuart/_0211_ ),
    .B1(\soc/simpleuart/_0212_ ),
    .Y(\soc/simpleuart/_0213_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0764_  (.A(\soc/simpleuart/_0210_ ),
    .B(\soc/simpleuart/_0213_ ),
    .Y(\soc/simpleuart/_0214_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0765_  (.A(\soc/simpleuart_reg_div_do[19] ),
    .B(\soc/simpleuart/send_divcnt[19] ),
    .Y(\soc/simpleuart/_0215_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0766_  (.A(\soc/simpleuart_reg_div_do[18] ),
    .B(\soc/simpleuart/send_divcnt[18] ),
    .Y(\soc/simpleuart/_0216_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_0767_  (.A(\soc/simpleuart/_0214_ ),
    .B(\soc/simpleuart/_0215_ ),
    .C(\soc/simpleuart/_0216_ ),
    .Y(\soc/simpleuart/_0217_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0768_  (.A_N(\soc/simpleuart/send_divcnt[16] ),
    .B(\soc/simpleuart_reg_div_do[16] ),
    .Y(\soc/simpleuart/_0218_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0769_  (.A(\soc/simpleuart_reg_div_do[20] ),
    .B(\soc/simpleuart/send_divcnt[20] ),
    .X(\soc/simpleuart/_0219_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0770_  (.A(\soc/simpleuart_reg_div_do[23] ),
    .Y(\soc/simpleuart/_0220_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0771_  (.A(\soc/simpleuart/_0220_ ),
    .B(\soc/simpleuart/send_divcnt[23] ),
    .Y(\soc/simpleuart/_0221_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0772_  (.A_N(\soc/simpleuart/send_divcnt[23] ),
    .B(\soc/simpleuart_reg_div_do[23] ),
    .Y(\soc/simpleuart/_0222_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0774_  (.A(\soc/simpleuart_reg_div_do[22] ),
    .B(\soc/simpleuart/send_divcnt[22] ),
    .Y(\soc/simpleuart/_0224_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_0775_  (.A(\soc/simpleuart/_0221_ ),
    .B(\soc/simpleuart/_0222_ ),
    .C(\soc/simpleuart/_0224_ ),
    .Y(\soc/simpleuart/_0225_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0776_  (.A(\soc/simpleuart_reg_div_do[21] ),
    .B(\soc/simpleuart/send_divcnt[21] ),
    .X(\soc/simpleuart/_0226_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0777_  (.A(\soc/simpleuart/_0219_ ),
    .B(\soc/simpleuart/_0225_ ),
    .C(\soc/simpleuart/_0226_ ),
    .Y(\soc/simpleuart/_0227_ ));
 sky130_fd_sc_hd__inv_2 \soc/simpleuart/_0778_  (.A(\soc/simpleuart_reg_div_do[16] ),
    .Y(\soc/simpleuart/_0228_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0779_  (.A(\soc/simpleuart_reg_div_do[17] ),
    .B(\soc/simpleuart/send_divcnt[17] ),
    .X(\soc/simpleuart/_0229_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0780_  (.A1(\soc/simpleuart/_0228_ ),
    .A2(\soc/simpleuart/send_divcnt[16] ),
    .B1(\soc/simpleuart/_0229_ ),
    .Y(\soc/simpleuart/_0230_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_0781_  (.A(\soc/simpleuart/_0218_ ),
    .B(\soc/simpleuart/_0227_ ),
    .C(\soc/simpleuart/_0230_ ),
    .Y(\soc/simpleuart/_0231_ ));
 sky130_fd_sc_hd__nor4_2 \soc/simpleuart/_0782_  (.A(\soc/simpleuart/_0191_ ),
    .B(\soc/simpleuart/_0204_ ),
    .C(\soc/simpleuart/_0217_ ),
    .D(\soc/simpleuart/_0231_ ),
    .Y(\soc/simpleuart/_0232_ ));
 sky130_fd_sc_hd__inv_2 \soc/simpleuart/_0783_  (.A(\soc/simpleuart_reg_div_do[21] ),
    .Y(\soc/simpleuart/_0233_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0784_  (.A_N(\soc/simpleuart/send_divcnt[20] ),
    .B(\soc/simpleuart_reg_div_do[20] ),
    .Y(\soc/simpleuart/_0234_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0785_  (.A(\soc/simpleuart/_0233_ ),
    .B(\soc/simpleuart/send_divcnt[21] ),
    .C(\soc/simpleuart/_0234_ ),
    .X(\soc/simpleuart/_0235_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/simpleuart/_0786_  (.A_N(\soc/simpleuart/send_divcnt[22] ),
    .B(\soc/simpleuart/_0221_ ),
    .C(\soc/simpleuart_reg_div_do[22] ),
    .Y(\soc/simpleuart/_0236_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0787_  (.A(\soc/simpleuart/_0215_ ),
    .B(\soc/simpleuart/_0216_ ),
    .Y(\soc/simpleuart/_0237_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0788_  (.A(\soc/simpleuart_reg_div_do[17] ),
    .Y(\soc/simpleuart/_0238_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0789_  (.A(\soc/simpleuart/_0238_ ),
    .B(\soc/simpleuart/send_divcnt[17] ),
    .C(\soc/simpleuart/_0218_ ),
    .X(\soc/simpleuart/_0239_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0790_  (.A(\soc/simpleuart/_0237_ ),
    .B(\soc/simpleuart/_0239_ ),
    .Y(\soc/simpleuart/_0240_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0791_  (.A(\soc/simpleuart/send_divcnt[19] ),
    .Y(\soc/simpleuart/_0241_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0792_  (.A(\soc/simpleuart_reg_div_do[18] ),
    .Y(\soc/simpleuart/_0242_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0793_  (.A(\soc/simpleuart/_0242_ ),
    .B(\soc/simpleuart/send_divcnt[18] ),
    .Y(\soc/simpleuart/_0243_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0794_  (.A(\soc/simpleuart_reg_div_do[19] ),
    .B(\soc/simpleuart/_0241_ ),
    .C(\soc/simpleuart/_0243_ ),
    .X(\soc/simpleuart/_0244_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0795_  (.A1(\soc/simpleuart/_0240_ ),
    .A2(\soc/simpleuart/_0244_ ),
    .B1(\soc/simpleuart/_0227_ ),
    .Y(\soc/simpleuart/_0245_ ));
 sky130_fd_sc_hd__o2111a_1 \soc/simpleuart/_0796_  (.A1(\soc/simpleuart/_0225_ ),
    .A2(\soc/simpleuart/_0235_ ),
    .B1(\soc/simpleuart/_0236_ ),
    .C1(\soc/simpleuart/_0245_ ),
    .D1(\soc/simpleuart/_0222_ ),
    .X(\soc/simpleuart/_0246_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0797_  (.A1(\soc/simpleuart/_0202_ ),
    .A2(\soc/simpleuart/_0199_ ),
    .B1(\soc/simpleuart/_0200_ ),
    .Y(\soc/simpleuart/_0247_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0798_  (.A(\soc/simpleuart/_0197_ ),
    .B(\soc/simpleuart/_0247_ ),
    .Y(\soc/simpleuart/_0248_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_0799_  (.A(\soc/simpleuart/_0193_ ),
    .B(\soc/simpleuart/send_divcnt[27] ),
    .C(\soc/simpleuart/_0194_ ),
    .X(\soc/simpleuart/_0249_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/simpleuart/_0800_  (.A1(\soc/simpleuart/_0204_ ),
    .A2(\soc/simpleuart/_0246_ ),
    .B1(\soc/simpleuart/_0248_ ),
    .C1(\soc/simpleuart/_0249_ ),
    .Y(\soc/simpleuart/_0250_ ));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 \soc/simpleuart/_0801_  (.A(\soc/simpleuart/_0214_ ),
    .SLEEP_B(\soc/simpleuart/_0250_ ),
    .X(\soc/simpleuart/_0251_ ));
 sky130_fd_sc_hd__nor2_2 \soc/simpleuart/_0802_  (.A(\soc/simpleuart/send_bitcnt[3] ),
    .B(\soc/simpleuart/_0133_ ),
    .Y(\soc/simpleuart/_0252_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_0803_  (.A(\soc/simpleuart/send_divcnt[30] ),
    .B(\soc/simpleuart/_0207_ ),
    .C_N(\soc/simpleuart_reg_div_do[30] ),
    .Y(\soc/simpleuart/_0253_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0804_  (.A(\soc/simpleuart/_0252_ ),
    .B(\soc/simpleuart/_0206_ ),
    .C(\soc/simpleuart/_0253_ ),
    .Y(\soc/simpleuart/_0254_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_0805_  (.A1(\soc/simpleuart/_0210_ ),
    .A2(\soc/simpleuart/_0212_ ),
    .B1(\soc/simpleuart/_0254_ ),
    .Y(\soc/simpleuart/_0255_ ));
 sky130_fd_sc_hd__nor3_4 \soc/simpleuart/_0806_  (.A(\soc/simpleuart/_0232_ ),
    .B(\soc/simpleuart/_0251_ ),
    .C(\soc/simpleuart/_0255_ ),
    .Y(\soc/simpleuart/_0256_ ));
 sky130_fd_sc_hd__and2_4 \soc/simpleuart/_0808_  (.A(\soc/_012_ ),
    .B(\soc/simpleuart/_0252_ ),
    .X(\soc/simpleuart/_0258_ ));
 sky130_fd_sc_hd__nor2_8 \soc/simpleuart/_0809_  (.A(\soc/simpleuart/_0256_ ),
    .B(\soc/simpleuart/_0258_ ),
    .Y(\soc/simpleuart/_0259_ ));
 sky130_fd_sc_hd__nand2_4 \soc/simpleuart/_0811_  (.A(\soc/simpleuart/send_dummy ),
    .B(\soc/simpleuart/_0252_ ),
    .Y(\soc/simpleuart/_0261_ ));
 sky130_fd_sc_hd__nand2_4 \soc/simpleuart/_0812_  (.A(_074_),
    .B(\soc/simpleuart/_0261_ ),
    .Y(\soc/simpleuart/_0262_ ));
 sky130_fd_sc_hd__a221o_1 \soc/simpleuart/_0813_  (.A1(\soc/simpleuart/send_pattern[1] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0259_ ),
    .B2(net14),
    .C1(\soc/simpleuart/_0262_ ),
    .X(\soc/simpleuart/_0024_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0814_  (.A(\soc/simpleuart/send_pattern[1] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0263_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0816_  (.A1(\soc/simpleuart/send_pattern[2] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0258_ ),
    .B2(net285),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0265_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0817_  (.A(\soc/simpleuart/_0263_ ),
    .B(\soc/simpleuart/_0265_ ),
    .Y(\soc/simpleuart/_0025_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0818_  (.A(\soc/simpleuart/send_pattern[2] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0266_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0819_  (.A1(\soc/simpleuart/send_pattern[3] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0258_ ),
    .B2(net279),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0267_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0820_  (.A(\soc/simpleuart/_0266_ ),
    .B(\soc/simpleuart/_0267_ ),
    .Y(\soc/simpleuart/_0026_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0821_  (.A(\soc/simpleuart/send_pattern[3] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0268_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0822_  (.A1(\soc/simpleuart/send_pattern[4] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0258_ ),
    .B2(net270),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0269_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0823_  (.A(\soc/simpleuart/_0268_ ),
    .B(\soc/simpleuart/_0269_ ),
    .Y(\soc/simpleuart/_0027_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0824_  (.A(\soc/simpleuart/send_pattern[4] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0270_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0825_  (.A1(\soc/simpleuart/send_pattern[5] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0258_ ),
    .B2(net267),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0271_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0826_  (.A(\soc/simpleuart/_0270_ ),
    .B(\soc/simpleuart/_0271_ ),
    .Y(\soc/simpleuart/_0028_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0827_  (.A(\soc/simpleuart/send_pattern[5] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0272_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0828_  (.A1(\soc/simpleuart/send_pattern[6] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0258_ ),
    .B2(net265),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0273_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0829_  (.A(\soc/simpleuart/_0272_ ),
    .B(\soc/simpleuart/_0273_ ),
    .Y(\soc/simpleuart/_0029_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0830_  (.A(\soc/simpleuart/send_pattern[6] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0274_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0831_  (.A1(\soc/simpleuart/send_pattern[7] ),
    .A2(\soc/simpleuart/_0256_ ),
    .B1(\soc/simpleuart/_0258_ ),
    .B2(net263),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0275_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0832_  (.A(\soc/simpleuart/_0274_ ),
    .B(\soc/simpleuart/_0275_ ),
    .Y(\soc/simpleuart/_0030_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/simpleuart/_0833_  (.A_N(\soc/simpleuart/_0258_ ),
    .B(\soc/simpleuart/_0256_ ),
    .C(\soc/simpleuart/send_pattern[8] ),
    .Y(\soc/simpleuart/_0276_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_0834_  (.A1(net255),
    .A2(\soc/simpleuart/_0258_ ),
    .B1(\soc/simpleuart/_0259_ ),
    .B2(\soc/simpleuart/send_pattern[7] ),
    .C1(\soc/simpleuart/_0262_ ),
    .Y(\soc/simpleuart/_0277_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0835_  (.A(\soc/simpleuart/_0276_ ),
    .B(\soc/simpleuart/_0277_ ),
    .Y(\soc/simpleuart/_0031_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0836_  (.A(\soc/simpleuart/send_pattern[8] ),
    .Y(\soc/simpleuart/_0278_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/simpleuart/_0837_  (.A1(net253),
    .A2(\soc/simpleuart/_0258_ ),
    .B1(\soc/simpleuart/_0262_ ),
    .C1(\soc/simpleuart/_0256_ ),
    .Y(\soc/simpleuart/_0279_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0838_  (.A1(\soc/simpleuart/_0278_ ),
    .A2(\soc/simpleuart/_0258_ ),
    .B1(\soc/simpleuart/_0279_ ),
    .Y(\soc/simpleuart/_0032_ ));
 sky130_fd_sc_hd__nand3_4 \soc/simpleuart/_0839_  (.A(_074_),
    .B(\soc/simpleuart/_0259_ ),
    .C(\soc/simpleuart/_0261_ ),
    .Y(\soc/simpleuart/_0280_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0841_  (.A(\soc/simpleuart/send_divcnt[0] ),
    .B(\soc/simpleuart/_0280_ ),
    .Y(\soc/simpleuart/_0042_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0842_  (.A(\soc/simpleuart/send_divcnt[0] ),
    .B(\soc/simpleuart/send_divcnt[1] ),
    .Y(\soc/simpleuart/_0282_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0843_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0282_ ),
    .Y(\soc/simpleuart/_0043_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0845_  (.A1(\soc/simpleuart/send_divcnt[0] ),
    .A2(\soc/simpleuart/send_divcnt[1] ),
    .B1(\soc/simpleuart/send_divcnt[2] ),
    .Y(\soc/simpleuart/_0284_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_0846_  (.A(\soc/simpleuart/send_divcnt[0] ),
    .B(\soc/simpleuart/send_divcnt[2] ),
    .C(\soc/simpleuart/send_divcnt[1] ),
    .X(\soc/simpleuart/_0285_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0847_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0284_ ),
    .C(\soc/simpleuart/_0285_ ),
    .Y(\soc/simpleuart/_0044_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0848_  (.A(\soc/simpleuart/send_divcnt[3] ),
    .B(\soc/simpleuart/_0285_ ),
    .Y(\soc/simpleuart/_0286_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_0849_  (.A(\soc/simpleuart/send_divcnt[0] ),
    .B(\soc/simpleuart/send_divcnt[3] ),
    .C(\soc/simpleuart/send_divcnt[2] ),
    .D(\soc/simpleuart/send_divcnt[1] ),
    .X(\soc/simpleuart/_0287_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0850_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0286_ ),
    .C(\soc/simpleuart/_0287_ ),
    .Y(\soc/simpleuart/_0045_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0851_  (.A(\soc/simpleuart/send_divcnt[4] ),
    .B(\soc/simpleuart/_0287_ ),
    .Y(\soc/simpleuart/_0288_ ));
 sky130_fd_sc_hd__and2_0 \soc/simpleuart/_0852_  (.A(\soc/simpleuart/send_divcnt[4] ),
    .B(\soc/simpleuart/_0287_ ),
    .X(\soc/simpleuart/_0289_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0853_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0288_ ),
    .C(\soc/simpleuart/_0289_ ),
    .Y(\soc/simpleuart/_0046_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0854_  (.A(\soc/simpleuart/send_divcnt[5] ),
    .B(\soc/simpleuart/_0289_ ),
    .Y(\soc/simpleuart/_0290_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0855_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0290_ ),
    .Y(\soc/simpleuart/_0047_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0856_  (.A1(\soc/simpleuart/send_divcnt[5] ),
    .A2(\soc/simpleuart/_0289_ ),
    .B1(\soc/simpleuart/send_divcnt[6] ),
    .Y(\soc/simpleuart/_0291_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_0857_  (.A(\soc/simpleuart/send_divcnt[6] ),
    .B(\soc/simpleuart/send_divcnt[5] ),
    .C(\soc/simpleuart/send_divcnt[4] ),
    .D(\soc/simpleuart/_0287_ ),
    .X(\soc/simpleuart/_0292_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0858_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0291_ ),
    .C(\soc/simpleuart/_0292_ ),
    .Y(\soc/simpleuart/_0048_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0859_  (.A(\soc/simpleuart/send_divcnt[7] ),
    .B(\soc/simpleuart/_0292_ ),
    .Y(\soc/simpleuart/_0293_ ));
 sky130_fd_sc_hd__and2_0 \soc/simpleuart/_0860_  (.A(\soc/simpleuart/send_divcnt[7] ),
    .B(\soc/simpleuart/_0292_ ),
    .X(\soc/simpleuart/_0294_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0861_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0293_ ),
    .C(\soc/simpleuart/_0294_ ),
    .Y(\soc/simpleuart/_0049_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0862_  (.A(\soc/simpleuart/send_divcnt[8] ),
    .B(\soc/simpleuart/_0294_ ),
    .Y(\soc/simpleuart/_0295_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0863_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0295_ ),
    .Y(\soc/simpleuart/_0050_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_0864_  (.A(\soc/simpleuart/send_divcnt[9] ),
    .B(\soc/simpleuart/send_divcnt[8] ),
    .C(\soc/simpleuart/send_divcnt[7] ),
    .D(\soc/simpleuart/_0292_ ),
    .X(\soc/simpleuart/_0296_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0865_  (.A1(\soc/simpleuart/send_divcnt[8] ),
    .A2(\soc/simpleuart/_0294_ ),
    .B1(\soc/simpleuart/send_divcnt[9] ),
    .Y(\soc/simpleuart/_0297_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0866_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0296_ ),
    .C(\soc/simpleuart/_0297_ ),
    .Y(\soc/simpleuart/_0051_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0867_  (.A(\soc/simpleuart/send_divcnt[10] ),
    .B(\soc/simpleuart/_0296_ ),
    .Y(\soc/simpleuart/_0298_ ));
 sky130_fd_sc_hd__and2_0 \soc/simpleuart/_0868_  (.A(\soc/simpleuart/send_divcnt[10] ),
    .B(\soc/simpleuart/_0296_ ),
    .X(\soc/simpleuart/_0299_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0869_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0298_ ),
    .C(\soc/simpleuart/_0299_ ),
    .Y(\soc/simpleuart/_0052_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0870_  (.A(\soc/simpleuart/send_divcnt[11] ),
    .B(\soc/simpleuart/_0299_ ),
    .Y(\soc/simpleuart/_0300_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0871_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0300_ ),
    .Y(\soc/simpleuart/_0053_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0872_  (.A1(\soc/simpleuart/send_divcnt[11] ),
    .A2(\soc/simpleuart/_0299_ ),
    .B1(\soc/simpleuart/send_divcnt[12] ),
    .Y(\soc/simpleuart/_0301_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_0873_  (.A(\soc/simpleuart/send_divcnt[12] ),
    .B(\soc/simpleuart/send_divcnt[11] ),
    .C(\soc/simpleuart/send_divcnt[10] ),
    .D(\soc/simpleuart/_0296_ ),
    .X(\soc/simpleuart/_0302_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0874_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0301_ ),
    .C(\soc/simpleuart/_0302_ ),
    .Y(\soc/simpleuart/_0054_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0875_  (.A(\soc/simpleuart/send_divcnt[13] ),
    .B(\soc/simpleuart/_0302_ ),
    .Y(\soc/simpleuart/_0303_ ));
 sky130_fd_sc_hd__and2_1 \soc/simpleuart/_0876_  (.A(\soc/simpleuart/send_divcnt[13] ),
    .B(\soc/simpleuart/_0302_ ),
    .X(\soc/simpleuart/_0304_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0877_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0303_ ),
    .C(\soc/simpleuart/_0304_ ),
    .Y(\soc/simpleuart/_0055_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0878_  (.A(\soc/simpleuart/send_divcnt[14] ),
    .B(\soc/simpleuart/_0304_ ),
    .Y(\soc/simpleuart/_0305_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0879_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0305_ ),
    .Y(\soc/simpleuart/_0056_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0881_  (.A1(\soc/simpleuart/send_divcnt[14] ),
    .A2(\soc/simpleuart/_0304_ ),
    .B1(\soc/simpleuart/send_divcnt[15] ),
    .Y(\soc/simpleuart/_0307_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_0882_  (.A(\soc/simpleuart/send_divcnt[15] ),
    .B(\soc/simpleuart/send_divcnt[14] ),
    .C(\soc/simpleuart/send_divcnt[13] ),
    .D(\soc/simpleuart/_0302_ ),
    .X(\soc/simpleuart/_0308_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0883_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0307_ ),
    .C(\soc/simpleuart/_0308_ ),
    .Y(\soc/simpleuart/_0057_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0884_  (.A(\soc/simpleuart/send_divcnt[16] ),
    .B(\soc/simpleuart/_0308_ ),
    .Y(\soc/simpleuart/_0309_ ));
 sky130_fd_sc_hd__and2_1 \soc/simpleuart/_0885_  (.A(\soc/simpleuart/send_divcnt[16] ),
    .B(\soc/simpleuart/_0308_ ),
    .X(\soc/simpleuart/_0310_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0886_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0309_ ),
    .C(\soc/simpleuart/_0310_ ),
    .Y(\soc/simpleuart/_0058_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0887_  (.A(\soc/simpleuart/send_divcnt[17] ),
    .B(\soc/simpleuart/_0310_ ),
    .Y(\soc/simpleuart/_0311_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0888_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0311_ ),
    .Y(\soc/simpleuart/_0059_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0889_  (.A1(\soc/simpleuart/send_divcnt[17] ),
    .A2(\soc/simpleuart/_0310_ ),
    .B1(\soc/simpleuart/send_divcnt[18] ),
    .Y(\soc/simpleuart/_0312_ ));
 sky130_fd_sc_hd__nand4_2 \soc/simpleuart/_0890_  (.A(\soc/simpleuart/send_divcnt[18] ),
    .B(\soc/simpleuart/send_divcnt[17] ),
    .C(\soc/simpleuart/send_divcnt[16] ),
    .D(\soc/simpleuart/_0308_ ),
    .Y(\soc/simpleuart/_0313_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_0891_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0312_ ),
    .C_N(\soc/simpleuart/_0313_ ),
    .Y(\soc/simpleuart/_0060_ ));
 sky130_fd_sc_hd__nor2_2 \soc/simpleuart/_0892_  (.A(\soc/simpleuart/_0241_ ),
    .B(\soc/simpleuart/_0313_ ),
    .Y(\soc/simpleuart/_0314_ ));
 sky130_fd_sc_hd__or2_0 \soc/simpleuart/_0893_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0314_ ),
    .X(\soc/simpleuart/_0315_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0894_  (.A1(\soc/simpleuart/_0241_ ),
    .A2(\soc/simpleuart/_0313_ ),
    .B1(\soc/simpleuart/_0315_ ),
    .Y(\soc/simpleuart/_0061_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0895_  (.A(\soc/simpleuart/send_divcnt[20] ),
    .B(\soc/simpleuart/_0314_ ),
    .Y(\soc/simpleuart/_0316_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0896_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0316_ ),
    .Y(\soc/simpleuart/_0062_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0897_  (.A(\soc/simpleuart/send_divcnt[20] ),
    .B(\soc/simpleuart/_0314_ ),
    .Y(\soc/simpleuart/_0317_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_0898_  (.A(\soc/simpleuart/send_divcnt[21] ),
    .B(\soc/simpleuart/_0317_ ),
    .X(\soc/simpleuart/_0318_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0899_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0318_ ),
    .Y(\soc/simpleuart/_0063_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_0900_  (.A(\soc/simpleuart/send_divcnt[22] ),
    .B(\soc/simpleuart/send_divcnt[21] ),
    .C(\soc/simpleuart/send_divcnt[20] ),
    .D(\soc/simpleuart/_0314_ ),
    .X(\soc/simpleuart/_0319_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_0901_  (.A1(\soc/simpleuart/send_divcnt[21] ),
    .A2(\soc/simpleuart/send_divcnt[20] ),
    .A3(\soc/simpleuart/_0314_ ),
    .B1(\soc/simpleuart/send_divcnt[22] ),
    .Y(\soc/simpleuart/_0320_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0902_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0319_ ),
    .C(\soc/simpleuart/_0320_ ),
    .Y(\soc/simpleuart/_0064_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/simpleuart/_0903_  (.A1(\soc/simpleuart/send_divcnt[23] ),
    .A2(\soc/simpleuart/_0319_ ),
    .B1_N(\soc/simpleuart/_0280_ ),
    .Y(\soc/simpleuart/_0321_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0904_  (.A1(\soc/simpleuart/send_divcnt[23] ),
    .A2(\soc/simpleuart/_0319_ ),
    .B1(\soc/simpleuart/_0321_ ),
    .Y(\soc/simpleuart/_0065_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_0905_  (.A(\soc/simpleuart/send_divcnt[24] ),
    .B(\soc/simpleuart/send_divcnt[23] ),
    .C(\soc/simpleuart/_0319_ ),
    .X(\soc/simpleuart/_0322_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0906_  (.A1(\soc/simpleuart/send_divcnt[23] ),
    .A2(\soc/simpleuart/_0319_ ),
    .B1(\soc/simpleuart/send_divcnt[24] ),
    .Y(\soc/simpleuart/_0323_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0907_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0322_ ),
    .C(\soc/simpleuart/_0323_ ),
    .Y(\soc/simpleuart/_0066_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_0908_  (.A(\soc/simpleuart/send_divcnt[25] ),
    .B(\soc/simpleuart/send_divcnt[24] ),
    .C(\soc/simpleuart/send_divcnt[23] ),
    .D(\soc/simpleuart/_0319_ ),
    .X(\soc/simpleuart/_0324_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0909_  (.A(\soc/simpleuart/send_divcnt[25] ),
    .B(\soc/simpleuart/_0322_ ),
    .Y(\soc/simpleuart/_0325_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0910_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0324_ ),
    .C(\soc/simpleuart/_0325_ ),
    .Y(\soc/simpleuart/_0067_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/simpleuart/_0911_  (.A1(\soc/simpleuart/send_divcnt[26] ),
    .A2(\soc/simpleuart/_0324_ ),
    .B1_N(\soc/simpleuart/_0280_ ),
    .Y(\soc/simpleuart/_0326_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0912_  (.A1(\soc/simpleuart/send_divcnt[26] ),
    .A2(\soc/simpleuart/_0324_ ),
    .B1(\soc/simpleuart/_0326_ ),
    .Y(\soc/simpleuart/_0068_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0913_  (.A1(\soc/simpleuart/send_divcnt[26] ),
    .A2(\soc/simpleuart/_0324_ ),
    .B1(\soc/simpleuart/send_divcnt[27] ),
    .Y(\soc/simpleuart/_0327_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_0914_  (.A(\soc/simpleuart/send_divcnt[27] ),
    .B(\soc/simpleuart/send_divcnt[26] ),
    .C(\soc/simpleuart/_0324_ ),
    .Y(\soc/simpleuart/_0328_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_0915_  (.A(\soc/simpleuart/_0327_ ),
    .B(\soc/simpleuart/_0280_ ),
    .C_N(\soc/simpleuart/_0328_ ),
    .Y(\soc/simpleuart/_0069_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0916_  (.A(\soc/simpleuart/_0211_ ),
    .B(\soc/simpleuart/_0328_ ),
    .Y(\soc/simpleuart/_0329_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_0917_  (.A1(\soc/simpleuart/send_divcnt[27] ),
    .A2(\soc/simpleuart/send_divcnt[26] ),
    .A3(\soc/simpleuart/_0324_ ),
    .B1(\soc/simpleuart/send_divcnt[28] ),
    .Y(\soc/simpleuart/_0330_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0918_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0329_ ),
    .C(\soc/simpleuart/_0330_ ),
    .Y(\soc/simpleuart/_0070_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/simpleuart/_0919_  (.A1(\soc/simpleuart/send_divcnt[29] ),
    .A2(\soc/simpleuart/_0329_ ),
    .B1_N(\soc/simpleuart/_0280_ ),
    .Y(\soc/simpleuart/_0331_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0920_  (.A1(\soc/simpleuart/send_divcnt[29] ),
    .A2(\soc/simpleuart/_0329_ ),
    .B1(\soc/simpleuart/_0331_ ),
    .Y(\soc/simpleuart/_0071_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_0921_  (.A(\soc/simpleuart/send_divcnt[30] ),
    .B(\soc/simpleuart/send_divcnt[29] ),
    .C(\soc/simpleuart/_0329_ ),
    .X(\soc/simpleuart/_0332_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0922_  (.A1(\soc/simpleuart/send_divcnt[29] ),
    .A2(\soc/simpleuart/_0329_ ),
    .B1(\soc/simpleuart/send_divcnt[30] ),
    .Y(\soc/simpleuart/_0333_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_0923_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0332_ ),
    .C(\soc/simpleuart/_0333_ ),
    .Y(\soc/simpleuart/_0072_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_0924_  (.A(\soc/simpleuart/send_divcnt[31] ),
    .B(\soc/simpleuart/_0332_ ),
    .Y(\soc/simpleuart/_0334_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0925_  (.A(\soc/simpleuart/_0280_ ),
    .B(\soc/simpleuart/_0334_ ),
    .Y(\soc/simpleuart/_0073_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0926_  (.A(\soc/simpleuart_reg_div_do[24] ),
    .B(net546),
    .Y(\soc/simpleuart/_0335_ ));
 sky130_fd_sc_hd__inv_2 \soc/simpleuart/_0927_  (.A(net546),
    .Y(\soc/simpleuart/_0336_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0929_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net185),
    .B1(_074_),
    .Y(\soc/simpleuart/_0338_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0930_  (.A(net547),
    .B(\soc/simpleuart/_0338_ ),
    .Y(\soc/simpleuart/_0000_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0931_  (.A(\soc/simpleuart_reg_div_do[25] ),
    .Y(\soc/simpleuart/_0339_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0934_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net182),
    .B1(_074_),
    .Y(\soc/simpleuart/_0342_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0935_  (.A1(\soc/simpleuart/_0339_ ),
    .A2(\soc/simpleuart/_0336_ ),
    .B1(\soc/simpleuart/_0342_ ),
    .Y(\soc/simpleuart/_0001_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0936_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net179),
    .B1(_074_),
    .Y(\soc/simpleuart/_0343_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0937_  (.A1(\soc/simpleuart/_0192_ ),
    .A2(\soc/simpleuart/_0336_ ),
    .B1(\soc/simpleuart/_0343_ ),
    .Y(\soc/simpleuart/_0002_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0938_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net176),
    .B1(_074_),
    .Y(\soc/simpleuart/_0344_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0939_  (.A1(\soc/simpleuart/_0193_ ),
    .A2(\soc/simpleuart/_0336_ ),
    .B1(\soc/simpleuart/_0344_ ),
    .Y(\soc/simpleuart/_0003_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0940_  (.A(\soc/simpleuart_reg_div_do[28] ),
    .Y(\soc/simpleuart/_0345_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0941_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net173),
    .B1(_074_),
    .Y(\soc/simpleuart/_0346_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0942_  (.A1(\soc/simpleuart/_0345_ ),
    .A2(\soc/simpleuart/_0336_ ),
    .B1(\soc/simpleuart/_0346_ ),
    .Y(\soc/simpleuart/_0004_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0943_  (.A(\soc/simpleuart_reg_div_do[29] ),
    .Y(\soc/simpleuart/_0347_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_0944_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net169),
    .B1(_074_),
    .Y(\soc/simpleuart/_0348_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0945_  (.A1(\soc/simpleuart/_0347_ ),
    .A2(\soc/simpleuart/_0336_ ),
    .B1(\soc/simpleuart/_0348_ ),
    .Y(\soc/simpleuart/_0005_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0946_  (.A(\soc/simpleuart_reg_div_do[30] ),
    .B(\soc/_011_ ),
    .Y(\soc/simpleuart/_0349_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0947_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net167),
    .B1(_074_),
    .Y(\soc/simpleuart/_0350_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0948_  (.A(\soc/simpleuart/_0349_ ),
    .B(\soc/simpleuart/_0350_ ),
    .Y(\soc/simpleuart/_0006_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0949_  (.A(\soc/simpleuart_reg_div_do[31] ),
    .B(\soc/_011_ ),
    .Y(\soc/simpleuart/_0351_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0950_  (.A1(\soc/simpleuart/_0336_ ),
    .A2(net165),
    .B1(_074_),
    .Y(\soc/simpleuart/_0352_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0951_  (.A(\soc/simpleuart/_0351_ ),
    .B(\soc/simpleuart/_0352_ ),
    .Y(\soc/simpleuart/_0007_ ));
 sky130_fd_sc_hd__clkinv_4 \soc/simpleuart/_0952_  (.A(\soc/_010_ ),
    .Y(\soc/simpleuart/_0353_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0954_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net212),
    .B1(_074_),
    .Y(\soc/simpleuart/_0355_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0955_  (.A1(\soc/simpleuart/_0228_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0355_ ),
    .Y(\soc/simpleuart/_0008_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0956_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net209),
    .B1(_074_),
    .Y(\soc/simpleuart/_0356_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0957_  (.A1(\soc/simpleuart/_0238_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0356_ ),
    .Y(\soc/simpleuart/_0009_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0958_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net206),
    .B1(_074_),
    .Y(\soc/simpleuart/_0357_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0959_  (.A1(\soc/simpleuart/_0242_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0357_ ),
    .Y(\soc/simpleuart/_0010_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0960_  (.A(\soc/simpleuart_reg_div_do[19] ),
    .Y(\soc/simpleuart/_0358_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0961_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net202),
    .B1(_074_),
    .Y(\soc/simpleuart/_0359_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0962_  (.A1(\soc/simpleuart/_0358_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0359_ ),
    .Y(\soc/simpleuart/_0011_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0963_  (.A(\soc/simpleuart_reg_div_do[20] ),
    .Y(\soc/simpleuart/_0360_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0965_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net199),
    .B1(_074_),
    .Y(\soc/simpleuart/_0362_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0966_  (.A1(\soc/simpleuart/_0360_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0362_ ),
    .Y(\soc/simpleuart/_0012_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0967_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net195),
    .B1(_074_),
    .Y(\soc/simpleuart/_0363_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0968_  (.A1(\soc/simpleuart/_0233_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0363_ ),
    .Y(\soc/simpleuart/_0013_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0969_  (.A(\soc/simpleuart_reg_div_do[22] ),
    .B(\soc/_010_ ),
    .Y(\soc/simpleuart/_0364_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0970_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net192),
    .B1(_074_),
    .Y(\soc/simpleuart/_0365_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_0971_  (.A(\soc/simpleuart/_0364_ ),
    .B(\soc/simpleuart/_0365_ ),
    .Y(\soc/simpleuart/_0014_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0972_  (.A1(\soc/simpleuart/_0353_ ),
    .A2(net188),
    .B1(_074_),
    .Y(\soc/simpleuart/_0366_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0973_  (.A1(\soc/simpleuart/_0220_ ),
    .A2(\soc/simpleuart/_0353_ ),
    .B1(\soc/simpleuart/_0366_ ),
    .Y(\soc/simpleuart/_0015_ ));
 sky130_fd_sc_hd__clkinv_4 \soc/simpleuart/_0974_  (.A(\soc/_009_ ),
    .Y(\soc/simpleuart/_0367_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0976_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net245),
    .B1(_074_),
    .Y(\soc/simpleuart/_0369_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0977_  (.A1(\soc/simpleuart/_0165_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0369_ ),
    .Y(\soc/simpleuart/_0016_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0978_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net237),
    .B1(_074_),
    .Y(\soc/simpleuart/_0370_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0979_  (.A1(\soc/simpleuart/_0170_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0370_ ),
    .Y(\soc/simpleuart/_0017_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0980_  (.A(\soc/simpleuart_reg_div_do[10] ),
    .Y(\soc/simpleuart/_0371_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0981_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net235),
    .B1(_074_),
    .Y(\soc/simpleuart/_0372_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0982_  (.A1(\soc/simpleuart/_0371_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0372_ ),
    .Y(\soc/simpleuart/_0018_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0983_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net231),
    .B1(_074_),
    .Y(\soc/simpleuart/_0373_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0984_  (.A1(\soc/simpleuart/_0172_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0373_ ),
    .Y(\soc/simpleuart/_0019_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0985_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net227),
    .B1(_074_),
    .Y(\soc/simpleuart/_0374_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0986_  (.A1(\soc/simpleuart/_0177_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0374_ ),
    .Y(\soc/simpleuart/_0020_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0987_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net223),
    .B1(_074_),
    .Y(\soc/simpleuart/_0375_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0988_  (.A1(\soc/simpleuart/_0178_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0375_ ),
    .Y(\soc/simpleuart/_0021_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_0989_  (.A(\soc/simpleuart_reg_div_do[14] ),
    .Y(\soc/simpleuart/_0376_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0990_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net220),
    .B1(_074_),
    .Y(\soc/simpleuart/_0377_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0991_  (.A1(\soc/simpleuart/_0376_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0377_ ),
    .Y(\soc/simpleuart/_0022_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_0993_  (.A1(\soc/simpleuart/_0367_ ),
    .A2(net216),
    .B1(_074_),
    .Y(\soc/simpleuart/_0379_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0994_  (.A1(\soc/simpleuart/_0187_ ),
    .A2(\soc/simpleuart/_0367_ ),
    .B1(\soc/simpleuart/_0379_ ),
    .Y(\soc/simpleuart/_0023_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_0995_  (.A(\soc/simpleuart/send_bitcnt[0] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0380_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_0996_  (.A_N(\soc/simpleuart/send_bitcnt[0] ),
    .B(\soc/simpleuart/_0256_ ),
    .Y(\soc/simpleuart/_0381_ ));
 sky130_fd_sc_hd__inv_2 \soc/simpleuart/_0997_  (.A(_074_),
    .Y(\soc/simpleuart/_0382_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_0998_  (.A1(\soc/simpleuart/_0261_ ),
    .A2(\soc/simpleuart/_0380_ ),
    .A3(\soc/simpleuart/_0381_ ),
    .B1(\soc/simpleuart/_0382_ ),
    .Y(\soc/simpleuart/_0033_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_0999_  (.A1(\soc/simpleuart/_0259_ ),
    .A2(\soc/simpleuart/_0261_ ),
    .B1(\soc/simpleuart/send_bitcnt[0] ),
    .Y(\soc/simpleuart/_0383_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1000_  (.A1(\soc/simpleuart/send_bitcnt[1] ),
    .A2(\soc/simpleuart/_0383_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0384_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1001_  (.A1(\soc/simpleuart/send_bitcnt[1] ),
    .A2(\soc/simpleuart/_0383_ ),
    .B1(\soc/simpleuart/_0384_ ),
    .Y(\soc/simpleuart/_0034_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1002_  (.A1(\soc/simpleuart/send_bitcnt[1] ),
    .A2(\soc/simpleuart/send_bitcnt[0] ),
    .B1(\soc/simpleuart/send_bitcnt[2] ),
    .Y(\soc/simpleuart/_0385_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1003_  (.A(\soc/simpleuart/_0133_ ),
    .B(\soc/simpleuart/_0385_ ),
    .Y(\soc/simpleuart/_0386_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1004_  (.A(\soc/simpleuart/_0256_ ),
    .B(\soc/simpleuart/_0386_ ),
    .Y(\soc/simpleuart/_0387_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1005_  (.A(\soc/simpleuart/send_bitcnt[2] ),
    .B(\soc/simpleuart/_0259_ ),
    .Y(\soc/simpleuart/_0388_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1006_  (.A1(\soc/simpleuart/_0261_ ),
    .A2(\soc/simpleuart/_0387_ ),
    .A3(\soc/simpleuart/_0388_ ),
    .B1(\soc/simpleuart/_0382_ ),
    .Y(\soc/simpleuart/_0035_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1007_  (.A1(\soc/simpleuart/_0133_ ),
    .A2(\soc/simpleuart/_0259_ ),
    .B1(\soc/simpleuart/send_bitcnt[3] ),
    .Y(\soc/simpleuart/_0389_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1008_  (.A(\soc/simpleuart/_0259_ ),
    .B(\soc/simpleuart/_0261_ ),
    .Y(\soc/simpleuart/_0390_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1009_  (.A(\soc/simpleuart/_0252_ ),
    .B(\soc/simpleuart/_0390_ ),
    .Y(\soc/simpleuart/_0391_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1010_  (.A1(\soc/simpleuart/_0389_ ),
    .A2(\soc/simpleuart/_0391_ ),
    .B1(\soc/simpleuart/_0382_ ),
    .Y(\soc/simpleuart/_0036_ ));
 sky130_fd_sc_hd__or4_1 \soc/simpleuart/_1011_  (.A(\soc/simpleuart/send_dummy ),
    .B(\soc/_009_ ),
    .C(\soc/_008_ ),
    .D(\soc/_010_ ),
    .X(\soc/simpleuart/_0392_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1012_  (.A1(\soc/_011_ ),
    .A2(\soc/simpleuart/_0392_ ),
    .B1(\soc/simpleuart/_0261_ ),
    .Y(\soc/simpleuart/_0393_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1013_  (.A(_074_),
    .B(\soc/simpleuart/_0393_ ),
    .Y(\soc/simpleuart/_0037_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1014_  (.A(\soc/simpleuart/recv_state[0] ),
    .Y(\soc/simpleuart/_0394_ ));
 sky130_fd_sc_hd__or3_2 \soc/simpleuart/_1015_  (.A(\soc/simpleuart/recv_state[1] ),
    .B(\soc/simpleuart/recv_state[2] ),
    .C(\soc/simpleuart/recv_state[3] ),
    .X(\soc/simpleuart/_0395_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1016_  (.A(\soc/simpleuart/recv_state[0] ),
    .B(\soc/simpleuart/_0395_ ),
    .Y(\soc/simpleuart/_0396_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1017_  (.A(\soc/simpleuart/recv_divcnt[5] ),
    .Y(\soc/simpleuart/_0397_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1018_  (.A(\soc/simpleuart/_0152_ ),
    .B(\soc/simpleuart/recv_divcnt[4] ),
    .Y(\soc/simpleuart/_0398_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1019_  (.A(\soc/simpleuart/recv_divcnt[2] ),
    .Y(\soc/simpleuart/_0399_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1020_  (.A_N(\soc/simpleuart_reg_div_do[1] ),
    .B(\soc/simpleuart/recv_divcnt[1] ),
    .Y(\soc/simpleuart/_0400_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1021_  (.A_N(\soc/simpleuart_reg_div_do[0] ),
    .B(\soc/simpleuart/recv_divcnt[0] ),
    .Y(\soc/simpleuart/_0401_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_1022_  (.A(\soc/simpleuart_reg_div_do[1] ),
    .SLEEP(\soc/simpleuart/recv_divcnt[1] ),
    .X(\soc/simpleuart/_0402_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_1023_  (.A1(\soc/simpleuart/_0399_ ),
    .A2(\soc/simpleuart_reg_div_do[2] ),
    .B1(\soc/simpleuart/_0400_ ),
    .B2(\soc/simpleuart/_0401_ ),
    .C1(\soc/simpleuart/_0402_ ),
    .Y(\soc/simpleuart/_0403_ ));
 sky130_fd_sc_hd__a22o_1 \soc/simpleuart/_1024_  (.A1(\soc/simpleuart/recv_divcnt[3] ),
    .A2(\soc/simpleuart/_0150_ ),
    .B1(\soc/simpleuart/recv_divcnt[2] ),
    .B2(\soc/simpleuart/_0145_ ),
    .X(\soc/simpleuart/_0404_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_1025_  (.A1(\soc/simpleuart/_0152_ ),
    .A2(\soc/simpleuart/recv_divcnt[4] ),
    .B1(\soc/simpleuart/recv_divcnt[3] ),
    .B2(\soc/simpleuart/_0150_ ),
    .Y(\soc/simpleuart/_0405_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/simpleuart/_1026_  (.A1(\soc/simpleuart/_0403_ ),
    .A2(\soc/simpleuart/_0404_ ),
    .B1_N(\soc/simpleuart/_0405_ ),
    .Y(\soc/simpleuart/_0406_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/simpleuart/_1027_  (.A1(\soc/simpleuart/_0397_ ),
    .A2(\soc/simpleuart_reg_div_do[5] ),
    .B1(\soc/simpleuart/_0398_ ),
    .B2(\soc/simpleuart/_0406_ ),
    .Y(\soc/simpleuart/_0407_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1028_  (.A(\soc/simpleuart/recv_divcnt[6] ),
    .Y(\soc/simpleuart/_0408_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/simpleuart/_1029_  (.A1(\soc/simpleuart/_0408_ ),
    .A2(\soc/simpleuart_reg_div_do[6] ),
    .B1(\soc/simpleuart/_0397_ ),
    .B2(\soc/simpleuart_reg_div_do[5] ),
    .Y(\soc/simpleuart/_0409_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1030_  (.A(\soc/simpleuart/_0408_ ),
    .B(\soc/simpleuart_reg_div_do[6] ),
    .Y(\soc/simpleuart/_0410_ ));
 sky130_fd_sc_hd__o221ai_4 \soc/simpleuart/_1031_  (.A1(\soc/simpleuart/recv_divcnt[7] ),
    .A2(\soc/simpleuart/_0159_ ),
    .B1(\soc/simpleuart/_0407_ ),
    .B2(\soc/simpleuart/_0409_ ),
    .C1(\soc/simpleuart/_0410_ ),
    .Y(\soc/simpleuart/_0411_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1032_  (.A_N(\soc/simpleuart/recv_divcnt[10] ),
    .B(\soc/simpleuart_reg_div_do[10] ),
    .Y(\soc/simpleuart/_0412_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1034_  (.A(\soc/simpleuart/recv_divcnt[11] ),
    .B(\soc/simpleuart_reg_div_do[11] ),
    .Y(\soc/simpleuart/_0414_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1035_  (.A(\soc/simpleuart/recv_divcnt[10] ),
    .B(\soc/simpleuart/_0371_ ),
    .Y(\soc/simpleuart/_0415_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_1036_  (.A(\soc/simpleuart/_0412_ ),
    .B(\soc/simpleuart/_0414_ ),
    .C(\soc/simpleuart/_0415_ ),
    .Y(\soc/simpleuart/_0416_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1038_  (.A(\soc/simpleuart/recv_divcnt[9] ),
    .B(\soc/simpleuart_reg_div_do[9] ),
    .X(\soc/simpleuart/_0418_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1039_  (.A(\soc/simpleuart/recv_divcnt[7] ),
    .Y(\soc/simpleuart/_0419_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1040_  (.A_N(\soc/simpleuart/recv_divcnt[8] ),
    .B(\soc/simpleuart_reg_div_do[8] ),
    .Y(\soc/simpleuart/_0420_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1041_  (.A1(\soc/simpleuart/_0419_ ),
    .A2(\soc/simpleuart_reg_div_do[7] ),
    .B1(\soc/simpleuart/_0420_ ),
    .Y(\soc/simpleuart/_0421_ ));
 sky130_fd_sc_hd__a2111oi_1 \soc/simpleuart/_1042_  (.A1(\soc/simpleuart/_0165_ ),
    .A2(\soc/simpleuart/recv_divcnt[8] ),
    .B1(\soc/simpleuart/_0416_ ),
    .C1(\soc/simpleuart/_0418_ ),
    .D1(\soc/simpleuart/_0421_ ),
    .Y(\soc/simpleuart/_0422_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1043_  (.A(\soc/simpleuart/recv_divcnt[9] ),
    .B(\soc/simpleuart/_0170_ ),
    .C(\soc/simpleuart/_0420_ ),
    .X(\soc/simpleuart/_0423_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1044_  (.A(\soc/simpleuart/recv_divcnt[11] ),
    .B(\soc/simpleuart/_0172_ ),
    .C(\soc/simpleuart/_0412_ ),
    .X(\soc/simpleuart/_0424_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1045_  (.A1(\soc/simpleuart/_0416_ ),
    .A2(\soc/simpleuart/_0423_ ),
    .B1(\soc/simpleuart/_0424_ ),
    .Y(\soc/simpleuart/_0425_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/simpleuart/_1046_  (.A1(\soc/simpleuart/_0411_ ),
    .A2(\soc/simpleuart/_0422_ ),
    .B1(\soc/simpleuart/_0425_ ),
    .Y(\soc/simpleuart/_0426_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1047_  (.A(\soc/simpleuart/recv_divcnt[15] ),
    .Y(\soc/simpleuart/_0427_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1048_  (.A(\soc/simpleuart/recv_divcnt[14] ),
    .B(\soc/simpleuart/_0376_ ),
    .Y(\soc/simpleuart/_0428_ ));
 sky130_fd_sc_hd__a22o_1 \soc/simpleuart/_1049_  (.A1(\soc/simpleuart/recv_divcnt[15] ),
    .A2(\soc/simpleuart/_0187_ ),
    .B1(\soc/simpleuart/recv_divcnt[14] ),
    .B2(\soc/simpleuart/_0376_ ),
    .X(\soc/simpleuart/_0429_ ));
 sky130_fd_sc_hd__a211o_1 \soc/simpleuart/_1050_  (.A1(\soc/simpleuart/_0427_ ),
    .A2(\soc/simpleuart_reg_div_do[15] ),
    .B1(\soc/simpleuart/_0428_ ),
    .C1(\soc/simpleuart/_0429_ ),
    .X(\soc/simpleuart/_0430_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1051_  (.A(\soc/simpleuart/recv_divcnt[13] ),
    .Y(\soc/simpleuart/_0431_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1052_  (.A(\soc/simpleuart/recv_divcnt[12] ),
    .Y(\soc/simpleuart/_0432_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_1053_  (.A1(\soc/simpleuart/_0431_ ),
    .A2(\soc/simpleuart_reg_div_do[13] ),
    .B1(\soc/simpleuart_reg_div_do[12] ),
    .B2(\soc/simpleuart/_0432_ ),
    .Y(\soc/simpleuart/_0433_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/simpleuart/_1054_  (.A1(\soc/simpleuart/recv_divcnt[13] ),
    .A2(\soc/simpleuart/_0178_ ),
    .B1(\soc/simpleuart/_0177_ ),
    .B2(\soc/simpleuart/recv_divcnt[12] ),
    .Y(\soc/simpleuart/_0434_ ));
 sky130_fd_sc_hd__nor4_2 \soc/simpleuart/_1055_  (.A(\soc/simpleuart/_0426_ ),
    .B(\soc/simpleuart/_0430_ ),
    .C(\soc/simpleuart/_0433_ ),
    .D(\soc/simpleuart/_0434_ ),
    .Y(\soc/simpleuart/_0435_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_1056_  (.A1(\soc/simpleuart/_0431_ ),
    .A2(\soc/simpleuart_reg_div_do[13] ),
    .B1(\soc/simpleuart/_0434_ ),
    .Y(\soc/simpleuart/_0436_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1057_  (.A(\soc/simpleuart/_0427_ ),
    .B(\soc/simpleuart_reg_div_do[15] ),
    .C(\soc/simpleuart/_0428_ ),
    .X(\soc/simpleuart/_0437_ ));
 sky130_fd_sc_hd__o21bai_2 \soc/simpleuart/_1058_  (.A1(\soc/simpleuart/_0430_ ),
    .A2(\soc/simpleuart/_0436_ ),
    .B1_N(\soc/simpleuart/_0437_ ),
    .Y(\soc/simpleuart/_0438_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1059_  (.A(net549),
    .B(\soc/simpleuart/_0238_ ),
    .Y(\soc/simpleuart/_0439_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1060_  (.A(net510),
    .B(\soc/simpleuart_reg_div_do[19] ),
    .X(\soc/simpleuart/_0440_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1061_  (.A(net538),
    .B(\soc/simpleuart_reg_div_do[18] ),
    .X(\soc/simpleuart/_0441_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/simpleuart/_1062_  (.A1(net549),
    .A2(\soc/simpleuart/_0238_ ),
    .B1(\soc/simpleuart/_0228_ ),
    .B2(\soc/simpleuart/recv_divcnt[16] ),
    .Y(\soc/simpleuart/_0442_ ));
 sky130_fd_sc_hd__a2111oi_0 \soc/simpleuart/_1063_  (.A1(\soc/simpleuart/_0228_ ),
    .A2(\soc/simpleuart/recv_divcnt[16] ),
    .B1(\soc/simpleuart/_0440_ ),
    .C1(\soc/simpleuart/_0441_ ),
    .D1(\soc/simpleuart/_0442_ ),
    .Y(\soc/simpleuart/_0443_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/simpleuart/_1064_  (.A1(\soc/simpleuart/_0435_ ),
    .A2(\soc/simpleuart/_0438_ ),
    .B1(net550),
    .C1(\soc/simpleuart/_0443_ ),
    .Y(\soc/simpleuart/_0444_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1065_  (.A(\soc/simpleuart/_0440_ ),
    .B(\soc/simpleuart/_0441_ ),
    .Y(\soc/simpleuart/_0445_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1066_  (.A(net510),
    .B(\soc/simpleuart/_0358_ ),
    .Y(\soc/simpleuart/_0446_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_1067_  (.A1(net510),
    .A2(\soc/simpleuart/_0358_ ),
    .B1(net538),
    .B2(\soc/simpleuart/_0242_ ),
    .Y(\soc/simpleuart/_0447_ ));
 sky130_fd_sc_hd__a32oi_2 \soc/simpleuart/_1068_  (.A1(\soc/simpleuart/_0445_ ),
    .A2(\soc/simpleuart/_0442_ ),
    .A3(net550),
    .B1(\soc/simpleuart/_0446_ ),
    .B2(\soc/simpleuart/_0447_ ),
    .Y(\soc/simpleuart/_0448_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1069_  (.A_N(\soc/simpleuart/recv_divcnt[26] ),
    .B(\soc/simpleuart_reg_div_do[26] ),
    .Y(\soc/simpleuart/_0449_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/simpleuart/_1070_  (.A1(\soc/simpleuart/recv_divcnt[27] ),
    .A2(\soc/simpleuart/_0193_ ),
    .B1(\soc/simpleuart/recv_divcnt[26] ),
    .B2(\soc/simpleuart/_0192_ ),
    .C1(\soc/simpleuart/recv_divcnt[25] ),
    .C2(\soc/simpleuart/_0339_ ),
    .Y(\soc/simpleuart/_0450_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/simpleuart/_1071_  (.A1(\soc/simpleuart/recv_divcnt[27] ),
    .A2(\soc/simpleuart/_0193_ ),
    .B1(\soc/simpleuart/_0449_ ),
    .C1(\soc/simpleuart/_0450_ ),
    .Y(\soc/simpleuart/_0451_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1072_  (.A(\soc/simpleuart/recv_divcnt[25] ),
    .B(\soc/simpleuart/_0339_ ),
    .Y(\soc/simpleuart/_0452_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1073_  (.A(\soc/simpleuart_reg_div_do[24] ),
    .B(\soc/simpleuart/recv_divcnt[24] ),
    .X(\soc/simpleuart/_0453_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1074_  (.A(\soc/simpleuart/_0451_ ),
    .B(\soc/simpleuart/_0452_ ),
    .C(\soc/simpleuart/_0453_ ),
    .Y(\soc/simpleuart/_0454_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1075_  (.A(\soc/simpleuart/recv_divcnt[30] ),
    .Y(\soc/simpleuart/_0455_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_1076_  (.A(\soc/simpleuart_reg_div_do[31] ),
    .SLEEP(\soc/simpleuart/recv_divcnt[31] ),
    .X(\soc/simpleuart/_0456_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1077_  (.A(\soc/simpleuart/recv_divcnt[29] ),
    .Y(\soc/simpleuart/_0457_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1078_  (.A_N(\soc/simpleuart_reg_div_do[31] ),
    .B(\soc/simpleuart/recv_divcnt[31] ),
    .Y(\soc/simpleuart/_0458_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/simpleuart/_1079_  (.A1(\soc/simpleuart/_0455_ ),
    .A2(\soc/simpleuart_reg_div_do[30] ),
    .B1(\soc/simpleuart/_0457_ ),
    .B2(\soc/simpleuart_reg_div_do[29] ),
    .C1(\soc/simpleuart/_0458_ ),
    .Y(\soc/simpleuart/_0459_ ));
 sky130_fd_sc_hd__a211o_1 \soc/simpleuart/_1080_  (.A1(\soc/simpleuart/_0455_ ),
    .A2(\soc/simpleuart_reg_div_do[30] ),
    .B1(\soc/simpleuart/_0456_ ),
    .C1(\soc/simpleuart/_0459_ ),
    .X(\soc/simpleuart/_0460_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1081_  (.A(\soc/simpleuart/recv_divcnt[28] ),
    .Y(\soc/simpleuart/_0461_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/simpleuart/_1082_  (.A1(\soc/simpleuart/_0457_ ),
    .A2(\soc/simpleuart_reg_div_do[29] ),
    .B1(\soc/simpleuart_reg_div_do[28] ),
    .B2(\soc/simpleuart/_0461_ ),
    .Y(\soc/simpleuart/_0462_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/simpleuart/_1083_  (.A1(\soc/simpleuart_reg_div_do[28] ),
    .A2(\soc/simpleuart/_0461_ ),
    .B1(\soc/simpleuart/_0462_ ),
    .Y(\soc/simpleuart/_0463_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/simpleuart/_1084_  (.A1(\soc/simpleuart/recv_divcnt[21] ),
    .A2(\soc/simpleuart/_0233_ ),
    .B1(\soc/simpleuart/_0360_ ),
    .B2(\soc/simpleuart/recv_divcnt[20] ),
    .Y(\soc/simpleuart/_0464_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1085_  (.A(\soc/simpleuart/recv_divcnt[21] ),
    .B(\soc/simpleuart/_0233_ ),
    .Y(\soc/simpleuart/_0465_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1086_  (.A(\soc/simpleuart/recv_divcnt[23] ),
    .B(\soc/simpleuart_reg_div_do[23] ),
    .Y(\soc/simpleuart/_0466_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1087_  (.A(\soc/simpleuart/recv_divcnt[22] ),
    .B(\soc/simpleuart_reg_div_do[22] ),
    .Y(\soc/simpleuart/_0467_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_1088_  (.A(\soc/simpleuart/_0465_ ),
    .B(\soc/simpleuart/_0466_ ),
    .C(\soc/simpleuart/_0467_ ),
    .Y(\soc/simpleuart/_0468_ ));
 sky130_fd_sc_hd__a21o_1 \soc/simpleuart/_1089_  (.A1(\soc/simpleuart/_0360_ ),
    .A2(\soc/simpleuart/recv_divcnt[20] ),
    .B1(\soc/simpleuart/_0468_ ),
    .X(\soc/simpleuart/_0469_ ));
 sky130_fd_sc_hd__nor4_1 \soc/simpleuart/_1090_  (.A(\soc/simpleuart/_0460_ ),
    .B(\soc/simpleuart/_0463_ ),
    .C(\soc/simpleuart/_0464_ ),
    .D(\soc/simpleuart/_0469_ ),
    .Y(\soc/simpleuart/_0470_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1091_  (.A(\soc/simpleuart/_0454_ ),
    .B(\soc/simpleuart/_0470_ ),
    .Y(\soc/simpleuart/_0471_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/simpleuart/_1092_  (.A1(\soc/simpleuart/_0444_ ),
    .A2(net551),
    .B1(\soc/simpleuart/_0471_ ),
    .Y(\soc/simpleuart/_0472_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1093_  (.A(\soc/simpleuart/recv_divcnt[23] ),
    .Y(\soc/simpleuart/_0473_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_1094_  (.A(\soc/simpleuart_reg_div_do[22] ),
    .SLEEP(\soc/simpleuart/recv_divcnt[22] ),
    .X(\soc/simpleuart/_0474_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1095_  (.A(\soc/simpleuart/_0473_ ),
    .B(\soc/simpleuart_reg_div_do[23] ),
    .C(\soc/simpleuart/_0474_ ),
    .X(\soc/simpleuart/_0475_ ));
 sky130_fd_sc_hd__a41o_1 \soc/simpleuart/_1096_  (.A1(\soc/simpleuart/_0465_ ),
    .A2(\soc/simpleuart/_0466_ ),
    .A3(\soc/simpleuart/_0467_ ),
    .A4(\soc/simpleuart/_0464_ ),
    .B1(\soc/simpleuart/_0475_ ),
    .X(\soc/simpleuart/_0476_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1097_  (.A(\soc/simpleuart/recv_divcnt[24] ),
    .Y(\soc/simpleuart/_0477_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1098_  (.A1(\soc/simpleuart_reg_div_do[24] ),
    .A2(\soc/simpleuart/_0477_ ),
    .B1(\soc/simpleuart/_0452_ ),
    .Y(\soc/simpleuart/_0478_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1099_  (.A(\soc/simpleuart/recv_divcnt[27] ),
    .B(\soc/simpleuart/_0193_ ),
    .C(\soc/simpleuart/_0449_ ),
    .X(\soc/simpleuart/_0479_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1100_  (.A1(\soc/simpleuart/_0451_ ),
    .A2(\soc/simpleuart/_0478_ ),
    .B1(\soc/simpleuart/_0479_ ),
    .Y(\soc/simpleuart/_0480_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1101_  (.A1(\soc/simpleuart/_0454_ ),
    .A2(\soc/simpleuart/_0476_ ),
    .B1(\soc/simpleuart/_0480_ ),
    .Y(\soc/simpleuart/_0481_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1102_  (.A(\soc/simpleuart/_0460_ ),
    .B(\soc/simpleuart/_0463_ ),
    .C(\soc/simpleuart/_0481_ ),
    .Y(\soc/simpleuart/_0482_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1103_  (.A1(\soc/simpleuart/_0455_ ),
    .A2(\soc/simpleuart_reg_div_do[30] ),
    .A3(\soc/simpleuart/_0458_ ),
    .B1(\soc/simpleuart/_0456_ ),
    .Y(\soc/simpleuart/_0483_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_1104_  (.A1(\soc/simpleuart/_0460_ ),
    .A2(\soc/simpleuart/_0462_ ),
    .B1(\soc/simpleuart/_0483_ ),
    .Y(\soc/simpleuart/_0484_ ));
 sky130_fd_sc_hd__nor3_4 \soc/simpleuart/_1105_  (.A(net552),
    .B(\soc/simpleuart/_0482_ ),
    .C(\soc/simpleuart/_0484_ ),
    .Y(\soc/simpleuart/_0485_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_1106_  (.A(\soc/simpleuart/recv_state[3] ),
    .SLEEP(\soc/simpleuart/recv_state[2] ),
    .X(\soc/simpleuart/_0486_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1107_  (.A(\soc/simpleuart/recv_state[1] ),
    .B(\soc/simpleuart/_0486_ ),
    .Y(\soc/simpleuart/_0487_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1108_  (.A(\soc/simpleuart/recv_state[0] ),
    .B(\soc/simpleuart/_0485_ ),
    .C(\soc/simpleuart/_0487_ ),
    .Y(\soc/simpleuart/_0488_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1109_  (.A(\soc/simpleuart_reg_div_do[3] ),
    .B(\soc/simpleuart/_0399_ ),
    .Y(\soc/simpleuart/_0489_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_1110_  (.A(\soc/simpleuart/recv_divcnt[0] ),
    .SLEEP(\soc/simpleuart_reg_div_do[1] ),
    .X(\soc/simpleuart/_0490_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1111_  (.A(\soc/simpleuart/_0145_ ),
    .B(\soc/simpleuart/recv_divcnt[1] ),
    .C(\soc/simpleuart/_0490_ ),
    .X(\soc/simpleuart/_0491_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1112_  (.A(\soc/simpleuart_reg_div_do[3] ),
    .B(\soc/simpleuart/_0399_ ),
    .Y(\soc/simpleuart/_0492_ ));
 sky130_fd_sc_hd__o221ai_2 \soc/simpleuart/_1113_  (.A1(\soc/simpleuart/_0152_ ),
    .A2(\soc/simpleuart/recv_divcnt[3] ),
    .B1(\soc/simpleuart/_0489_ ),
    .B2(\soc/simpleuart/_0491_ ),
    .C1(\soc/simpleuart/_0492_ ),
    .Y(\soc/simpleuart/_0493_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1114_  (.A(\soc/simpleuart/_0143_ ),
    .B(\soc/simpleuart/recv_divcnt[4] ),
    .Y(\soc/simpleuart/_0494_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1115_  (.A(\soc/simpleuart/_0152_ ),
    .B(\soc/simpleuart/recv_divcnt[3] ),
    .Y(\soc/simpleuart/_0495_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_1116_  (.A1(\soc/simpleuart/_0156_ ),
    .A2(\soc/simpleuart/recv_divcnt[5] ),
    .B1(\soc/simpleuart/_0143_ ),
    .B2(\soc/simpleuart/recv_divcnt[4] ),
    .Y(\soc/simpleuart/_0496_ ));
 sky130_fd_sc_hd__a31oi_2 \soc/simpleuart/_1117_  (.A1(\soc/simpleuart/_0493_ ),
    .A2(\soc/simpleuart/_0494_ ),
    .A3(\soc/simpleuart/_0495_ ),
    .B1(\soc/simpleuart/_0496_ ),
    .Y(\soc/simpleuart/_0497_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_1118_  (.A1(\soc/simpleuart_reg_div_do[7] ),
    .A2(\soc/simpleuart/_0408_ ),
    .B1(\soc/simpleuart_reg_div_do[6] ),
    .B2(\soc/simpleuart/_0397_ ),
    .Y(\soc/simpleuart/_0498_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/simpleuart/_1119_  (.A1(\soc/simpleuart_reg_div_do[8] ),
    .A2(\soc/simpleuart/_0419_ ),
    .B1(\soc/simpleuart_reg_div_do[7] ),
    .B2(\soc/simpleuart/_0408_ ),
    .Y(\soc/simpleuart/_0499_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_1120_  (.A1(\soc/simpleuart/_0497_ ),
    .A2(\soc/simpleuart/_0498_ ),
    .B1(\soc/simpleuart/_0499_ ),
    .Y(\soc/simpleuart/_0500_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1121_  (.A_N(\soc/simpleuart/recv_divcnt[10] ),
    .B(\soc/simpleuart_reg_div_do[11] ),
    .Y(\soc/simpleuart/_0501_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1122_  (.A(\soc/simpleuart/_0172_ ),
    .B(\soc/simpleuart/recv_divcnt[10] ),
    .Y(\soc/simpleuart/_0502_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1123_  (.A(\soc/simpleuart_reg_div_do[12] ),
    .B(\soc/simpleuart/recv_divcnt[11] ),
    .Y(\soc/simpleuart/_0503_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_1124_  (.A(\soc/simpleuart/_0501_ ),
    .B(\soc/simpleuart/_0502_ ),
    .C(\soc/simpleuart/_0503_ ),
    .Y(\soc/simpleuart/_0504_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1125_  (.A_N(\soc/simpleuart/recv_divcnt[8] ),
    .B(\soc/simpleuart_reg_div_do[9] ),
    .Y(\soc/simpleuart/_0505_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/simpleuart/_1126_  (.A1(\soc/simpleuart/_0371_ ),
    .A2(\soc/simpleuart/recv_divcnt[9] ),
    .B1(\soc/simpleuart_reg_div_do[8] ),
    .B2(\soc/simpleuart/_0419_ ),
    .Y(\soc/simpleuart/_0506_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/simpleuart/_1127_  (.A1(\soc/simpleuart/_0371_ ),
    .A2(\soc/simpleuart/recv_divcnt[9] ),
    .B1(\soc/simpleuart/_0170_ ),
    .B2(\soc/simpleuart/recv_divcnt[8] ),
    .C1(\soc/simpleuart/_0506_ ),
    .Y(\soc/simpleuart/_0507_ ));
 sky130_fd_sc_hd__and3b_1 \soc/simpleuart/_1128_  (.A_N(\soc/simpleuart/_0504_ ),
    .B(\soc/simpleuart/_0505_ ),
    .C(\soc/simpleuart/_0507_ ),
    .X(\soc/simpleuart/_0508_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1129_  (.A(\soc/simpleuart/_0371_ ),
    .B(\soc/simpleuart/recv_divcnt[9] ),
    .C(\soc/simpleuart/_0505_ ),
    .X(\soc/simpleuart/_0509_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1130_  (.A(\soc/simpleuart/_0177_ ),
    .B(\soc/simpleuart/recv_divcnt[11] ),
    .C(\soc/simpleuart/_0501_ ),
    .X(\soc/simpleuart/_0510_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_1131_  (.A1(\soc/simpleuart/_0504_ ),
    .A2(\soc/simpleuart/_0509_ ),
    .B1(\soc/simpleuart/_0510_ ),
    .Y(\soc/simpleuart/_0511_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/simpleuart/_1132_  (.A1(\soc/simpleuart/_0500_ ),
    .A2(\soc/simpleuart/_0508_ ),
    .B1(\soc/simpleuart/_0511_ ),
    .Y(\soc/simpleuart/_0512_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1133_  (.A(\soc/simpleuart/_0187_ ),
    .B(\soc/simpleuart/recv_divcnt[14] ),
    .Y(\soc/simpleuart/_0513_ ));
 sky130_fd_sc_hd__a22o_1 \soc/simpleuart/_1134_  (.A1(\soc/simpleuart/_0228_ ),
    .A2(\soc/simpleuart/recv_divcnt[15] ),
    .B1(\soc/simpleuart/_0187_ ),
    .B2(\soc/simpleuart/recv_divcnt[14] ),
    .X(\soc/simpleuart/_0514_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/simpleuart/_1135_  (.A1(\soc/simpleuart_reg_div_do[16] ),
    .A2(\soc/simpleuart/_0427_ ),
    .B1(\soc/simpleuart/_0513_ ),
    .C1(\soc/simpleuart/_0514_ ),
    .Y(\soc/simpleuart/_0515_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/simpleuart/_1136_  (.A1(\soc/simpleuart_reg_div_do[14] ),
    .A2(\soc/simpleuart/_0431_ ),
    .B1(\soc/simpleuart_reg_div_do[13] ),
    .B2(\soc/simpleuart/_0432_ ),
    .Y(\soc/simpleuart/_0516_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/simpleuart/_1137_  (.A1(\soc/simpleuart/_0376_ ),
    .A2(\soc/simpleuart/recv_divcnt[13] ),
    .B1(\soc/simpleuart/_0178_ ),
    .B2(\soc/simpleuart/recv_divcnt[12] ),
    .Y(\soc/simpleuart/_0517_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_1138_  (.A(\soc/simpleuart/_0515_ ),
    .B(\soc/simpleuart/_0516_ ),
    .C(\soc/simpleuart/_0517_ ),
    .Y(\soc/simpleuart/_0518_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1139_  (.A1(\soc/simpleuart/_0376_ ),
    .A2(\soc/simpleuart/recv_divcnt[13] ),
    .B1(\soc/simpleuart/_0516_ ),
    .Y(\soc/simpleuart/_0519_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1140_  (.A(\soc/simpleuart_reg_div_do[16] ),
    .B(\soc/simpleuart/_0427_ ),
    .C(\soc/simpleuart/_0513_ ),
    .X(\soc/simpleuart/_0520_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1141_  (.A1(\soc/simpleuart/_0515_ ),
    .A2(\soc/simpleuart/_0519_ ),
    .B1(\soc/simpleuart/_0520_ ),
    .Y(\soc/simpleuart/_0521_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/simpleuart/_1142_  (.A1(\soc/simpleuart/_0512_ ),
    .A2(\soc/simpleuart/_0518_ ),
    .B1(\soc/simpleuart/_0521_ ),
    .Y(\soc/simpleuart/_0522_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1143_  (.A(\soc/simpleuart/recv_divcnt[21] ),
    .Y(\soc/simpleuart/_0523_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1144_  (.A(\soc/simpleuart/_0220_ ),
    .B(\soc/simpleuart/recv_divcnt[22] ),
    .Y(\soc/simpleuart/_0524_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/simpleuart/_1145_  (.A(\soc/simpleuart/recv_divcnt[22] ),
    .SLEEP(\soc/simpleuart_reg_div_do[23] ),
    .X(\soc/simpleuart/_0525_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1146_  (.A(\soc/simpleuart_reg_div_do[24] ),
    .B(\soc/simpleuart/recv_divcnt[23] ),
    .X(\soc/simpleuart/_0526_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1147_  (.A(\soc/simpleuart/_0524_ ),
    .B(\soc/simpleuart/_0525_ ),
    .C(\soc/simpleuart/_0526_ ),
    .Y(\soc/simpleuart/_0527_ ));
 sky130_fd_sc_hd__o21a_1 \soc/simpleuart/_1148_  (.A1(\soc/simpleuart_reg_div_do[22] ),
    .A2(\soc/simpleuart/_0523_ ),
    .B1(\soc/simpleuart/_0527_ ),
    .X(\soc/simpleuart/_0528_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \soc/simpleuart/_1149_  (.A1_N(\soc/simpleuart/recv_divcnt[20] ),
    .A2_N(\soc/simpleuart/_0233_ ),
    .B1(\soc/simpleuart/_0523_ ),
    .B2(\soc/simpleuart_reg_div_do[22] ),
    .Y(\soc/simpleuart/_0529_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1150_  (.A(\soc/simpleuart/_0233_ ),
    .B(\soc/simpleuart/recv_divcnt[20] ),
    .Y(\soc/simpleuart/_0530_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1151_  (.A_N(\soc/simpleuart/recv_divcnt[16] ),
    .B(\soc/simpleuart_reg_div_do[17] ),
    .Y(\soc/simpleuart/_0531_ ));
 sky130_fd_sc_hd__nand4_1 \soc/simpleuart/_1152_  (.A(\soc/simpleuart/_0528_ ),
    .B(\soc/simpleuart/_0529_ ),
    .C(\soc/simpleuart/_0530_ ),
    .D(\soc/simpleuart/_0531_ ),
    .Y(\soc/simpleuart/_0532_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1153_  (.A(\soc/simpleuart_reg_div_do[19] ),
    .B(net538),
    .Y(\soc/simpleuart/_0533_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1154_  (.A(\soc/simpleuart_reg_div_do[20] ),
    .B(net510),
    .Y(\soc/simpleuart/_0534_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1155_  (.A(\soc/simpleuart_reg_div_do[18] ),
    .B(net549),
    .Y(\soc/simpleuart/_0535_ ));
 sky130_fd_sc_hd__nand3_1 \soc/simpleuart/_1156_  (.A(\soc/simpleuart/_0533_ ),
    .B(\soc/simpleuart/_0534_ ),
    .C(\soc/simpleuart/_0535_ ),
    .Y(\soc/simpleuart/_0536_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/simpleuart/_1157_  (.A1(\soc/simpleuart/_0238_ ),
    .A2(\soc/simpleuart/recv_divcnt[16] ),
    .B1(\soc/simpleuart/_0532_ ),
    .C1(\soc/simpleuart/_0536_ ),
    .Y(\soc/simpleuart/_0537_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1158_  (.A(\soc/simpleuart_reg_div_do[24] ),
    .B(\soc/simpleuart/_0473_ ),
    .C(\soc/simpleuart/_0524_ ),
    .X(\soc/simpleuart/_0538_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1159_  (.A1(\soc/simpleuart_reg_div_do[22] ),
    .A2(\soc/simpleuart/_0523_ ),
    .B1(\soc/simpleuart/_0527_ ),
    .Y(\soc/simpleuart/_0539_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1160_  (.A(\soc/simpleuart/_0533_ ),
    .B(\soc/simpleuart/_0534_ ),
    .Y(\soc/simpleuart/_0540_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1161_  (.A(\soc/simpleuart/_0242_ ),
    .B(net549),
    .C(\soc/simpleuart/_0531_ ),
    .X(\soc/simpleuart/_0541_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1162_  (.A_N(net538),
    .B(\soc/simpleuart_reg_div_do[19] ),
    .Y(\soc/simpleuart/_0542_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1163_  (.A(\soc/simpleuart/_0360_ ),
    .B(net510),
    .C(\soc/simpleuart/_0542_ ),
    .X(\soc/simpleuart/_0543_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1164_  (.A1(\soc/simpleuart/_0540_ ),
    .A2(\soc/simpleuart/_0541_ ),
    .B1(\soc/simpleuart/_0543_ ),
    .Y(\soc/simpleuart/_0544_ ));
 sky130_fd_sc_hd__nand4_1 \soc/simpleuart/_1165_  (.A(\soc/simpleuart/_0528_ ),
    .B(\soc/simpleuart/_0529_ ),
    .C(\soc/simpleuart/_0530_ ),
    .D(\soc/simpleuart/_0544_ ),
    .Y(\soc/simpleuart/_0545_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/simpleuart/_1166_  (.A1(\soc/simpleuart/_0539_ ),
    .A2(\soc/simpleuart/_0529_ ),
    .B1(\soc/simpleuart/_0545_ ),
    .Y(\soc/simpleuart/_0546_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/simpleuart/_1167_  (.A1(\soc/simpleuart/_0522_ ),
    .A2(\soc/simpleuart/_0537_ ),
    .B1(\soc/simpleuart/_0538_ ),
    .C1(\soc/simpleuart/_0546_ ),
    .Y(\soc/simpleuart/_0547_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1168_  (.A(\soc/simpleuart/_0192_ ),
    .B(\soc/simpleuart/recv_divcnt[25] ),
    .Y(\soc/simpleuart/_0548_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1169_  (.A(\soc/simpleuart_reg_div_do[27] ),
    .B(\soc/simpleuart/recv_divcnt[26] ),
    .Y(\soc/simpleuart/_0549_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1170_  (.A(\soc/simpleuart_reg_div_do[28] ),
    .B(\soc/simpleuart/recv_divcnt[27] ),
    .Y(\soc/simpleuart/_0550_ ));
 sky130_fd_sc_hd__o22ai_2 \soc/simpleuart/_1171_  (.A1(\soc/simpleuart/_0192_ ),
    .A2(\soc/simpleuart/recv_divcnt[25] ),
    .B1(\soc/simpleuart/_0339_ ),
    .B2(\soc/simpleuart/recv_divcnt[24] ),
    .Y(\soc/simpleuart/_0551_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1172_  (.A1(\soc/simpleuart/_0339_ ),
    .A2(\soc/simpleuart/recv_divcnt[24] ),
    .B1(\soc/simpleuart/_0551_ ),
    .Y(\soc/simpleuart/_0552_ ));
 sky130_fd_sc_hd__nand4_2 \soc/simpleuart/_1173_  (.A(\soc/simpleuart/_0548_ ),
    .B(\soc/simpleuart/_0549_ ),
    .C(\soc/simpleuart/_0550_ ),
    .D(\soc/simpleuart/_0552_ ),
    .Y(\soc/simpleuart/_0553_ ));
 sky130_fd_sc_hd__nand4_2 \soc/simpleuart/_1174_  (.A(\soc/simpleuart/_0548_ ),
    .B(\soc/simpleuart/_0549_ ),
    .C(\soc/simpleuart/_0550_ ),
    .D(\soc/simpleuart/_0551_ ),
    .Y(\soc/simpleuart/_0554_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1175_  (.A_N(\soc/simpleuart/recv_divcnt[26] ),
    .B(\soc/simpleuart_reg_div_do[27] ),
    .Y(\soc/simpleuart/_0555_ ));
 sky130_fd_sc_hd__maj3_1 \soc/simpleuart/_1176_  (.A(\soc/simpleuart/_0345_ ),
    .B(\soc/simpleuart/recv_divcnt[27] ),
    .C(\soc/simpleuart/_0555_ ),
    .X(\soc/simpleuart/_0556_ ));
 sky130_fd_sc_hd__o211ai_4 \soc/simpleuart/_1177_  (.A1(\soc/simpleuart/_0547_ ),
    .A2(\soc/simpleuart/_0553_ ),
    .B1(\soc/simpleuart/_0554_ ),
    .C1(\soc/simpleuart/_0556_ ),
    .Y(\soc/simpleuart/_0557_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/simpleuart/_1178_  (.A1(\soc/simpleuart_reg_div_do[30] ),
    .A2(\soc/simpleuart/_0457_ ),
    .B1(\soc/simpleuart_reg_div_do[29] ),
    .B2(\soc/simpleuart/_0461_ ),
    .Y(\soc/simpleuart/_0558_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1179_  (.A(\soc/simpleuart_reg_div_do[30] ),
    .B(\soc/simpleuart/_0457_ ),
    .Y(\soc/simpleuart/_0559_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1180_  (.A1(\soc/simpleuart/_0347_ ),
    .A2(\soc/simpleuart/recv_divcnt[28] ),
    .B1(\soc/simpleuart/_0559_ ),
    .Y(\soc/simpleuart/_0560_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \soc/simpleuart/_1181_  (.A1_N(\soc/simpleuart_reg_div_do[31] ),
    .A2_N(\soc/simpleuart/_0455_ ),
    .B1(\soc/simpleuart/_0558_ ),
    .B2(\soc/simpleuart/_0559_ ),
    .Y(\soc/simpleuart/_0561_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/simpleuart/_1182_  (.A1(\soc/simpleuart/_0557_ ),
    .A2(\soc/simpleuart/_0558_ ),
    .A3(\soc/simpleuart/_0560_ ),
    .B1(\soc/simpleuart/_0561_ ),
    .Y(\soc/simpleuart/_0562_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/simpleuart/_1183_  (.A1(\soc/simpleuart_reg_div_do[31] ),
    .A2(\soc/simpleuart/_0455_ ),
    .B1(\soc/simpleuart/recv_state[0] ),
    .Y(\soc/simpleuart/_0563_ ));
 sky130_fd_sc_hd__nor2_4 \soc/simpleuart/_1184_  (.A(\soc/simpleuart/recv_state[0] ),
    .B(\soc/simpleuart/_0487_ ),
    .Y(\soc/simpleuart/_0564_ ));
 sky130_fd_sc_hd__nor2b_2 \soc/simpleuart/_1185_  (.A(\soc/simpleuart/_0564_ ),
    .B_N(\soc/simpleuart/_0395_ ),
    .Y(\soc/simpleuart/_0565_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1186_  (.A(\soc/simpleuart/_0565_ ),
    .Y(\soc/simpleuart/_0566_ ));
 sky130_fd_sc_hd__o32ai_4 \soc/simpleuart/_1187_  (.A1(\soc/simpleuart/_0395_ ),
    .A2(\soc/simpleuart/_0562_ ),
    .A3(\soc/simpleuart/_0563_ ),
    .B1(\soc/simpleuart/_0566_ ),
    .B2(net553),
    .Y(\soc/simpleuart/_0567_ ));
 sky130_fd_sc_hd__a211o_1 \soc/simpleuart/_1188_  (.A1(net1),
    .A2(\soc/simpleuart/_0396_ ),
    .B1(\soc/simpleuart/_0488_ ),
    .C1(\soc/simpleuart/_0567_ ),
    .X(\soc/simpleuart/_0568_ ));
 sky130_fd_sc_hd__nor3_2 \soc/simpleuart/_1189_  (.A(\soc/simpleuart/_0394_ ),
    .B(\soc/simpleuart/_0567_ ),
    .C(\soc/simpleuart/_0488_ ),
    .Y(\soc/simpleuart/_0569_ ));
 sky130_fd_sc_hd__a2111oi_0 \soc/simpleuart/_1190_  (.A1(\soc/simpleuart/_0394_ ),
    .A2(\soc/simpleuart/_0568_ ),
    .B1(\soc/simpleuart/_0569_ ),
    .C1(\soc/simpleuart/_0382_ ),
    .D1(\soc/simpleuart/_0564_ ),
    .Y(\soc/simpleuart/_0038_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1191_  (.A(\soc/simpleuart/recv_state[0] ),
    .B(\soc/simpleuart/_0486_ ),
    .Y(\soc/simpleuart/_0570_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1192_  (.A(\soc/simpleuart/_0570_ ),
    .B(\soc/simpleuart/_0568_ ),
    .C_N(\soc/simpleuart/recv_state[1] ),
    .Y(\soc/simpleuart/_0571_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1193_  (.A1(\soc/simpleuart/recv_state[1] ),
    .A2(\soc/simpleuart/_0569_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0572_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1194_  (.A(\soc/simpleuart/_0571_ ),
    .B(\soc/simpleuart/_0572_ ),
    .Y(\soc/simpleuart/_0039_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_1195_  (.A(\soc/simpleuart/recv_state[1] ),
    .B(\soc/simpleuart/recv_state[2] ),
    .C(\soc/simpleuart/_0569_ ),
    .X(\soc/simpleuart/_0573_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1196_  (.A1(\soc/simpleuart/recv_state[1] ),
    .A2(\soc/simpleuart/_0569_ ),
    .B1(\soc/simpleuart/recv_state[2] ),
    .Y(\soc/simpleuart/_0574_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1197_  (.A(\soc/simpleuart/_0382_ ),
    .B(\soc/simpleuart/_0573_ ),
    .C(\soc/simpleuart/_0574_ ),
    .Y(\soc/simpleuart/_0040_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_1198_  (.A(\soc/simpleuart/recv_state[1] ),
    .B(\soc/simpleuart/recv_state[2] ),
    .C(\soc/simpleuart/recv_state[3] ),
    .D(\soc/simpleuart/_0569_ ),
    .X(\soc/simpleuart/_0575_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1199_  (.A1(\soc/simpleuart/_0565_ ),
    .A2(\soc/simpleuart/_0568_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0576_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1200_  (.A1(\soc/simpleuart/recv_state[1] ),
    .A2(\soc/simpleuart/recv_state[2] ),
    .A3(\soc/simpleuart/_0569_ ),
    .B1(\soc/simpleuart/recv_state[3] ),
    .Y(\soc/simpleuart/_0577_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1201_  (.A(\soc/simpleuart/_0575_ ),
    .B(\soc/simpleuart/_0576_ ),
    .C(\soc/simpleuart/_0577_ ),
    .Y(\soc/simpleuart/_0041_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1202_  (.A(\soc/simpleuart/recv_pattern[0] ),
    .Y(\soc/simpleuart/_0578_ ));
 sky130_fd_sc_hd__nand2_8 \soc/simpleuart/_1203_  (.A(\soc/simpleuart/_0485_ ),
    .B(\soc/simpleuart/_0565_ ),
    .Y(\soc/simpleuart/_0579_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1205_  (.A1(\soc/simpleuart/recv_pattern[1] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0581_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1206_  (.A1(\soc/simpleuart/_0578_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0581_ ),
    .Y(\soc/simpleuart/_0074_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1207_  (.A(\soc/simpleuart/recv_pattern[1] ),
    .Y(\soc/simpleuart/_0582_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1208_  (.A1(\soc/simpleuart/recv_pattern[2] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0583_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1209_  (.A1(\soc/simpleuart/_0582_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0583_ ),
    .Y(\soc/simpleuart/_0075_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1210_  (.A(\soc/simpleuart/recv_pattern[2] ),
    .Y(\soc/simpleuart/_0584_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1211_  (.A1(\soc/simpleuart/recv_pattern[3] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0585_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1212_  (.A1(\soc/simpleuart/_0584_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0585_ ),
    .Y(\soc/simpleuart/_0076_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1213_  (.A(\soc/simpleuart/recv_pattern[3] ),
    .Y(\soc/simpleuart/_0586_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1214_  (.A1(\soc/simpleuart/recv_pattern[4] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0587_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1215_  (.A1(\soc/simpleuart/_0586_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0587_ ),
    .Y(\soc/simpleuart/_0077_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1216_  (.A(\soc/simpleuart/recv_pattern[4] ),
    .Y(\soc/simpleuart/_0588_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1217_  (.A1(\soc/simpleuart/recv_pattern[5] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0589_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1218_  (.A1(\soc/simpleuart/_0588_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0589_ ),
    .Y(\soc/simpleuart/_0078_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1219_  (.A(\soc/simpleuart/recv_pattern[5] ),
    .Y(\soc/simpleuart/_0590_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1220_  (.A1(\soc/simpleuart/recv_pattern[6] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0591_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1221_  (.A1(\soc/simpleuart/_0590_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0591_ ),
    .Y(\soc/simpleuart/_0079_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1222_  (.A(\soc/simpleuart/recv_pattern[6] ),
    .Y(\soc/simpleuart/_0592_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1223_  (.A1(\soc/simpleuart/recv_pattern[7] ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0593_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1224_  (.A1(\soc/simpleuart/_0592_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0593_ ),
    .Y(\soc/simpleuart/_0080_ ));
 sky130_fd_sc_hd__inv_1 \soc/simpleuart/_1225_  (.A(\soc/simpleuart/recv_pattern[7] ),
    .Y(\soc/simpleuart/_0594_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1226_  (.A1(net1),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0595_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1227_  (.A1(\soc/simpleuart/_0594_ ),
    .A2(\soc/simpleuart/_0579_ ),
    .B1(\soc/simpleuart/_0595_ ),
    .Y(\soc/simpleuart/_0081_ ));
 sky130_fd_sc_hd__nand2_8 \soc/simpleuart/_1228_  (.A(\soc/simpleuart/_0485_ ),
    .B(\soc/simpleuart/_0564_ ),
    .Y(\soc/simpleuart/_0596_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1231_  (.A1(\soc/simpleuart/recv_pattern[0] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0599_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1232_  (.A1(\soc/simpleuart/_0134_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0599_ ),
    .Y(\soc/simpleuart/_0082_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1233_  (.A1(\soc/simpleuart/recv_pattern[1] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0600_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1234_  (.A1(\soc/simpleuart/_0136_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0600_ ),
    .Y(\soc/simpleuart/_0083_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1235_  (.A1(\soc/simpleuart/recv_pattern[2] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0601_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1236_  (.A1(\soc/simpleuart/_0137_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0601_ ),
    .Y(\soc/simpleuart/_0084_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1237_  (.A1(\soc/simpleuart/recv_pattern[3] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0602_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1238_  (.A1(\soc/simpleuart/_0138_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0602_ ),
    .Y(\soc/simpleuart/_0085_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1239_  (.A1(\soc/simpleuart/recv_pattern[4] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0603_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1240_  (.A1(\soc/simpleuart/_0139_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0603_ ),
    .Y(\soc/simpleuart/_0086_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1241_  (.A1(\soc/simpleuart/recv_pattern[5] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0604_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1242_  (.A1(\soc/simpleuart/_0140_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0604_ ),
    .Y(\soc/simpleuart/_0087_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1243_  (.A1(\soc/simpleuart/recv_pattern[6] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0605_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1244_  (.A1(\soc/simpleuart/_0141_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0605_ ),
    .Y(\soc/simpleuart/_0088_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1245_  (.A1(\soc/simpleuart/recv_pattern[7] ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(_074_),
    .Y(\soc/simpleuart/_0606_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1246_  (.A1(\soc/simpleuart/_0142_ ),
    .A2(\soc/simpleuart/_0596_ ),
    .B1(\soc/simpleuart/_0606_ ),
    .Y(\soc/simpleuart/_0089_ ));
 sky130_fd_sc_hd__o21ai_4 \soc/simpleuart/_1247_  (.A1(\soc/simpleuart/_0564_ ),
    .A2(net554),
    .B1(_074_),
    .Y(\soc/simpleuart/_0607_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1249_  (.A(\soc/simpleuart/recv_divcnt[0] ),
    .B(net62),
    .Y(\soc/simpleuart/_0090_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1250_  (.A(\soc/simpleuart/recv_divcnt[1] ),
    .B(\soc/simpleuart/recv_divcnt[0] ),
    .Y(\soc/simpleuart/_0609_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1251_  (.A(net62),
    .B(\soc/simpleuart/_0609_ ),
    .Y(\soc/simpleuart/_0091_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_1253_  (.A(\soc/simpleuart/recv_divcnt[2] ),
    .B(\soc/simpleuart/recv_divcnt[1] ),
    .C(\soc/simpleuart/recv_divcnt[0] ),
    .X(\soc/simpleuart/_0611_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1254_  (.A1(\soc/simpleuart/recv_divcnt[1] ),
    .A2(\soc/simpleuart/recv_divcnt[0] ),
    .B1(\soc/simpleuart/recv_divcnt[2] ),
    .Y(\soc/simpleuart/_0612_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1255_  (.A(net62),
    .B(\soc/simpleuart/_0611_ ),
    .C(\soc/simpleuart/_0612_ ),
    .Y(\soc/simpleuart/_0092_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_1256_  (.A(\soc/simpleuart/recv_divcnt[3] ),
    .B(\soc/simpleuart/recv_divcnt[2] ),
    .C(\soc/simpleuart/recv_divcnt[1] ),
    .D(\soc/simpleuart/recv_divcnt[0] ),
    .X(\soc/simpleuart/_0613_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1257_  (.A(\soc/simpleuart/recv_divcnt[3] ),
    .B(\soc/simpleuart/_0611_ ),
    .Y(\soc/simpleuart/_0614_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1258_  (.A(net62),
    .B(\soc/simpleuart/_0613_ ),
    .C(\soc/simpleuart/_0614_ ),
    .Y(\soc/simpleuart/_0093_ ));
 sky130_fd_sc_hd__and2_1 \soc/simpleuart/_1259_  (.A(\soc/simpleuart/recv_divcnt[4] ),
    .B(\soc/simpleuart/_0613_ ),
    .X(\soc/simpleuart/_0615_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1260_  (.A(\soc/simpleuart/recv_divcnt[4] ),
    .B(\soc/simpleuart/_0613_ ),
    .Y(\soc/simpleuart/_0616_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1261_  (.A(net62),
    .B(\soc/simpleuart/_0615_ ),
    .C(\soc/simpleuart/_0616_ ),
    .Y(\soc/simpleuart/_0094_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1262_  (.A(\soc/simpleuart/recv_divcnt[5] ),
    .B(\soc/simpleuart/_0615_ ),
    .Y(\soc/simpleuart/_0617_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1263_  (.A(net62),
    .B(\soc/simpleuart/_0617_ ),
    .Y(\soc/simpleuart/_0095_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_1265_  (.A(\soc/simpleuart/recv_divcnt[6] ),
    .B(\soc/simpleuart/recv_divcnt[5] ),
    .C(\soc/simpleuart/_0615_ ),
    .X(\soc/simpleuart/_0619_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1266_  (.A1(\soc/simpleuart/recv_divcnt[5] ),
    .A2(\soc/simpleuart/_0615_ ),
    .B1(\soc/simpleuart/recv_divcnt[6] ),
    .Y(\soc/simpleuart/_0620_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1267_  (.A(net62),
    .B(\soc/simpleuart/_0619_ ),
    .C(\soc/simpleuart/_0620_ ),
    .Y(\soc/simpleuart/_0096_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_1268_  (.A(\soc/simpleuart/recv_divcnt[7] ),
    .B(\soc/simpleuart/recv_divcnt[6] ),
    .C(\soc/simpleuart/recv_divcnt[5] ),
    .D(\soc/simpleuart/_0615_ ),
    .X(\soc/simpleuart/_0621_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1269_  (.A(\soc/simpleuart/recv_divcnt[7] ),
    .B(\soc/simpleuart/_0619_ ),
    .Y(\soc/simpleuart/_0622_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1270_  (.A(net62),
    .B(\soc/simpleuart/_0621_ ),
    .C(\soc/simpleuart/_0622_ ),
    .Y(\soc/simpleuart/_0097_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1271_  (.A(\soc/simpleuart/recv_divcnt[8] ),
    .B(\soc/simpleuart/_0621_ ),
    .Y(\soc/simpleuart/_0623_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1272_  (.A(\soc/simpleuart/recv_divcnt[8] ),
    .B(\soc/simpleuart/_0621_ ),
    .Y(\soc/simpleuart/_0624_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1273_  (.A(\soc/simpleuart/_0623_ ),
    .B(net62),
    .C_N(\soc/simpleuart/_0624_ ),
    .Y(\soc/simpleuart/_0098_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1274_  (.A(\soc/simpleuart/recv_divcnt[9] ),
    .B(\soc/simpleuart/_0624_ ),
    .X(\soc/simpleuart/_0625_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1275_  (.A(net62),
    .B(\soc/simpleuart/_0625_ ),
    .Y(\soc/simpleuart/_0099_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_1276_  (.A(\soc/simpleuart/recv_divcnt[10] ),
    .B(\soc/simpleuart/recv_divcnt[9] ),
    .C(\soc/simpleuart/recv_divcnt[8] ),
    .D(\soc/simpleuart/_0621_ ),
    .X(\soc/simpleuart/_0626_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1277_  (.A1(\soc/simpleuart/recv_divcnt[9] ),
    .A2(\soc/simpleuart/recv_divcnt[8] ),
    .A3(\soc/simpleuart/_0621_ ),
    .B1(\soc/simpleuart/recv_divcnt[10] ),
    .Y(\soc/simpleuart/_0627_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1278_  (.A(net62),
    .B(\soc/simpleuart/_0626_ ),
    .C(\soc/simpleuart/_0627_ ),
    .Y(\soc/simpleuart/_0100_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1279_  (.A(\soc/simpleuart/recv_divcnt[11] ),
    .B(\soc/simpleuart/_0626_ ),
    .Y(\soc/simpleuart/_0628_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1280_  (.A(\soc/simpleuart/recv_divcnt[11] ),
    .B(\soc/simpleuart/_0626_ ),
    .Y(\soc/simpleuart/_0629_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1281_  (.A(\soc/simpleuart/_0628_ ),
    .B(net62),
    .C_N(\soc/simpleuart/_0629_ ),
    .Y(\soc/simpleuart/_0101_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1282_  (.A(\soc/simpleuart/_0432_ ),
    .B(\soc/simpleuart/_0629_ ),
    .Y(\soc/simpleuart/_0630_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1283_  (.A(net62),
    .B(\soc/simpleuart/_0630_ ),
    .Y(\soc/simpleuart/_0102_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_1284_  (.A(\soc/simpleuart/recv_divcnt[13] ),
    .B(\soc/simpleuart/recv_divcnt[12] ),
    .C(\soc/simpleuart/recv_divcnt[11] ),
    .D(\soc/simpleuart/_0626_ ),
    .X(\soc/simpleuart/_0631_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1285_  (.A1(\soc/simpleuart/recv_divcnt[12] ),
    .A2(\soc/simpleuart/recv_divcnt[11] ),
    .A3(\soc/simpleuart/_0626_ ),
    .B1(\soc/simpleuart/recv_divcnt[13] ),
    .Y(\soc/simpleuart/_0632_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1286_  (.A(net62),
    .B(\soc/simpleuart/_0631_ ),
    .C(\soc/simpleuart/_0632_ ),
    .Y(\soc/simpleuart/_0103_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1287_  (.A(\soc/simpleuart/recv_divcnt[14] ),
    .B(\soc/simpleuart/_0631_ ),
    .Y(\soc/simpleuart/_0633_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1288_  (.A(\soc/simpleuart/recv_divcnt[14] ),
    .B(\soc/simpleuart/_0631_ ),
    .Y(\soc/simpleuart/_0634_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1289_  (.A(\soc/simpleuart/_0633_ ),
    .B(net62),
    .C_N(\soc/simpleuart/_0634_ ),
    .Y(\soc/simpleuart/_0104_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1290_  (.A(\soc/simpleuart/_0427_ ),
    .B(\soc/simpleuart/_0634_ ),
    .Y(\soc/simpleuart/_0635_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1291_  (.A(net62),
    .B(\soc/simpleuart/_0635_ ),
    .Y(\soc/simpleuart/_0105_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_1292_  (.A(\soc/simpleuart/recv_divcnt[16] ),
    .B(\soc/simpleuart/recv_divcnt[15] ),
    .C(\soc/simpleuart/recv_divcnt[14] ),
    .D(\soc/simpleuart/_0631_ ),
    .X(\soc/simpleuart/_0636_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1293_  (.A1(\soc/simpleuart/recv_divcnt[15] ),
    .A2(\soc/simpleuart/recv_divcnt[14] ),
    .A3(\soc/simpleuart/_0631_ ),
    .B1(\soc/simpleuart/recv_divcnt[16] ),
    .Y(\soc/simpleuart/_0637_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1294_  (.A(net62),
    .B(\soc/simpleuart/_0636_ ),
    .C(\soc/simpleuart/_0637_ ),
    .Y(\soc/simpleuart/_0106_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1295_  (.A(\soc/simpleuart/recv_divcnt[17] ),
    .B(\soc/simpleuart/_0636_ ),
    .Y(\soc/simpleuart/_0638_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1296_  (.A(\soc/simpleuart/recv_divcnt[17] ),
    .B(\soc/simpleuart/_0636_ ),
    .Y(\soc/simpleuart/_0639_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1297_  (.A(\soc/simpleuart/_0638_ ),
    .B(\soc/simpleuart/_0607_ ),
    .C_N(\soc/simpleuart/_0639_ ),
    .Y(\soc/simpleuart/_0107_ ));
 sky130_fd_sc_hd__xor2_1 \soc/simpleuart/_1298_  (.A(\soc/simpleuart/recv_divcnt[18] ),
    .B(\soc/simpleuart/_0639_ ),
    .X(\soc/simpleuart/_0640_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1299_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0640_ ),
    .Y(\soc/simpleuart/_0108_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_1300_  (.A(net510),
    .B(net538),
    .C(\soc/simpleuart/recv_divcnt[17] ),
    .D(\soc/simpleuart/_0636_ ),
    .X(\soc/simpleuart/_0641_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1301_  (.A1(\soc/simpleuart/recv_divcnt[18] ),
    .A2(\soc/simpleuart/recv_divcnt[17] ),
    .A3(\soc/simpleuart/_0636_ ),
    .B1(\soc/simpleuart/recv_divcnt[19] ),
    .Y(\soc/simpleuart/_0642_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1302_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0641_ ),
    .C(\soc/simpleuart/_0642_ ),
    .Y(\soc/simpleuart/_0109_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1303_  (.A(\soc/simpleuart/recv_divcnt[20] ),
    .B(net511),
    .Y(\soc/simpleuart/_0643_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1304_  (.A(\soc/simpleuart/recv_divcnt[20] ),
    .B(net511),
    .Y(\soc/simpleuart/_0644_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1305_  (.A(\soc/simpleuart/_0643_ ),
    .B(\soc/simpleuart/_0607_ ),
    .C_N(\soc/simpleuart/_0644_ ),
    .Y(\soc/simpleuart/_0110_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1306_  (.A(\soc/simpleuart/_0523_ ),
    .B(\soc/simpleuart/_0644_ ),
    .Y(\soc/simpleuart/_0645_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1307_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0645_ ),
    .Y(\soc/simpleuart/_0111_ ));
 sky130_fd_sc_hd__and4_1 \soc/simpleuart/_1308_  (.A(\soc/simpleuart/recv_divcnt[22] ),
    .B(net921),
    .C(net707),
    .D(net540),
    .X(\soc/simpleuart/_0646_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1309_  (.A1(net921),
    .A2(net707),
    .A3(net540),
    .B1(\soc/simpleuart/recv_divcnt[22] ),
    .Y(\soc/simpleuart/_0647_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1310_  (.A(net555),
    .B(net541),
    .C(net512),
    .Y(\soc/simpleuart/_0112_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1311_  (.A(\soc/simpleuart/recv_divcnt[23] ),
    .B(net541),
    .Y(\soc/simpleuart/_0648_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1312_  (.A(\soc/simpleuart/recv_divcnt[23] ),
    .B(net541),
    .Y(\soc/simpleuart/_0649_ ));
 sky130_fd_sc_hd__nor3b_1 \soc/simpleuart/_1313_  (.A(net542),
    .B(net555),
    .C_N(\soc/simpleuart/_0649_ ),
    .Y(\soc/simpleuart/_0113_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1314_  (.A(\soc/simpleuart/_0477_ ),
    .B(\soc/simpleuart/_0649_ ),
    .Y(\soc/simpleuart/_0650_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1315_  (.A(net555),
    .B(\soc/simpleuart/_0650_ ),
    .Y(\soc/simpleuart/_0114_ ));
 sky130_fd_sc_hd__and4_2 \soc/simpleuart/_1316_  (.A(\soc/simpleuart/recv_divcnt[25] ),
    .B(\soc/simpleuart/recv_divcnt[24] ),
    .C(\soc/simpleuart/recv_divcnt[23] ),
    .D(\soc/simpleuart/_0646_ ),
    .X(\soc/simpleuart/_0651_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/simpleuart/_1317_  (.A1(\soc/simpleuart/recv_divcnt[24] ),
    .A2(\soc/simpleuart/recv_divcnt[23] ),
    .A3(\soc/simpleuart/_0646_ ),
    .B1(\soc/simpleuart/recv_divcnt[25] ),
    .Y(\soc/simpleuart/_0652_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1318_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0651_ ),
    .C(\soc/simpleuart/_0652_ ),
    .Y(\soc/simpleuart/_0115_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1319_  (.A(\soc/simpleuart/recv_divcnt[26] ),
    .B(\soc/simpleuart/_0651_ ),
    .Y(\soc/simpleuart/_0653_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1320_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0653_ ),
    .Y(\soc/simpleuart/_0116_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_1321_  (.A(\soc/simpleuart/recv_divcnt[27] ),
    .B(\soc/simpleuart/recv_divcnt[26] ),
    .C(\soc/simpleuart/_0651_ ),
    .X(\soc/simpleuart/_0654_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1322_  (.A1(\soc/simpleuart/recv_divcnt[26] ),
    .A2(\soc/simpleuart/_0651_ ),
    .B1(\soc/simpleuart/recv_divcnt[27] ),
    .Y(\soc/simpleuart/_0655_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1323_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0654_ ),
    .C(\soc/simpleuart/_0655_ ),
    .Y(\soc/simpleuart/_0117_ ));
 sky130_fd_sc_hd__and2_1 \soc/simpleuart/_1324_  (.A(\soc/simpleuart/recv_divcnt[28] ),
    .B(\soc/simpleuart/_0654_ ),
    .X(\soc/simpleuart/_0656_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1325_  (.A(\soc/simpleuart/recv_divcnt[28] ),
    .B(\soc/simpleuart/_0654_ ),
    .Y(\soc/simpleuart/_0657_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1326_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0656_ ),
    .C(\soc/simpleuart/_0657_ ),
    .Y(\soc/simpleuart/_0118_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/simpleuart/_1327_  (.A1(\soc/simpleuart/recv_divcnt[29] ),
    .A2(\soc/simpleuart/_0656_ ),
    .B1_N(\soc/simpleuart/_0607_ ),
    .Y(\soc/simpleuart/_0658_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1328_  (.A1(\soc/simpleuart/recv_divcnt[29] ),
    .A2(\soc/simpleuart/_0656_ ),
    .B1(\soc/simpleuart/_0658_ ),
    .Y(\soc/simpleuart/_0119_ ));
 sky130_fd_sc_hd__and3_1 \soc/simpleuart/_1329_  (.A(\soc/simpleuart/recv_divcnt[30] ),
    .B(\soc/simpleuart/recv_divcnt[29] ),
    .C(\soc/simpleuart/_0656_ ),
    .X(\soc/simpleuart/_0659_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1330_  (.A1(\soc/simpleuart/recv_divcnt[29] ),
    .A2(\soc/simpleuart/_0656_ ),
    .B1(\soc/simpleuart/recv_divcnt[30] ),
    .Y(\soc/simpleuart/_0660_ ));
 sky130_fd_sc_hd__nor3_1 \soc/simpleuart/_1331_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0659_ ),
    .C(\soc/simpleuart/_0660_ ),
    .Y(\soc/simpleuart/_0120_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/simpleuart/_1332_  (.A(\soc/simpleuart/recv_divcnt[31] ),
    .B(\soc/simpleuart/_0659_ ),
    .Y(\soc/simpleuart/_0661_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1333_  (.A(\soc/simpleuart/_0607_ ),
    .B(\soc/simpleuart/_0661_ ),
    .Y(\soc/simpleuart/_0121_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1334_  (.A(\soc/_008_ ),
    .B(net285),
    .Y(\soc/simpleuart/_0662_ ));
 sky130_fd_sc_hd__inv_2 \soc/simpleuart/_1335_  (.A(\soc/_008_ ),
    .Y(\soc/simpleuart/_0663_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1337_  (.A1(\soc/simpleuart_reg_div_do[0] ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0382_ ),
    .Y(\soc/simpleuart/_0665_ ));
 sky130_fd_sc_hd__nand2_1 \soc/simpleuart/_1338_  (.A(\soc/simpleuart/_0662_ ),
    .B(\soc/simpleuart/_0665_ ),
    .Y(\soc/simpleuart/_0122_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1339_  (.A(\soc/simpleuart_reg_div_do[1] ),
    .B(\soc/_008_ ),
    .Y(\soc/simpleuart/_0666_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1340_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net279),
    .B1(_074_),
    .Y(\soc/simpleuart/_0667_ ));
 sky130_fd_sc_hd__nor2_1 \soc/simpleuart/_1341_  (.A(\soc/simpleuart/_0666_ ),
    .B(\soc/simpleuart/_0667_ ),
    .Y(\soc/simpleuart/_0123_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1342_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net270),
    .B1(_074_),
    .Y(\soc/simpleuart/_0668_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1343_  (.A1(\soc/simpleuart/_0145_ ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0668_ ),
    .Y(\soc/simpleuart/_0124_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1344_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net267),
    .B1(_074_),
    .Y(\soc/simpleuart/_0669_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1345_  (.A1(\soc/simpleuart/_0150_ ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0669_ ),
    .Y(\soc/simpleuart/_0125_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1346_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net265),
    .B1(_074_),
    .Y(\soc/simpleuart/_0670_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1347_  (.A1(\soc/simpleuart/_0152_ ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0670_ ),
    .Y(\soc/simpleuart/_0126_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1348_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net263),
    .B1(_074_),
    .Y(\soc/simpleuart/_0671_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1349_  (.A1(\soc/simpleuart/_0143_ ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0671_ ),
    .Y(\soc/simpleuart/_0127_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1350_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net255),
    .B1(_074_),
    .Y(\soc/simpleuart/_0672_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1351_  (.A1(\soc/simpleuart/_0156_ ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0672_ ),
    .Y(\soc/simpleuart/_0128_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/simpleuart/_1352_  (.A1(\soc/simpleuart/_0663_ ),
    .A2(net253),
    .B1(_074_),
    .Y(\soc/simpleuart/_0131_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1353_  (.A1(\soc/simpleuart/_0159_ ),
    .A2(\soc/simpleuart/_0663_ ),
    .B1(\soc/simpleuart/_0131_ ),
    .Y(\soc/simpleuart/_0129_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/simpleuart/_1354_  (.A_N(\soc/_002_ ),
    .B(\soc/simpleuart/recv_buf_valid ),
    .Y(\soc/simpleuart/_0132_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/simpleuart/_1355_  (.A1(\soc/simpleuart/_0596_ ),
    .A2(\soc/simpleuart/_0132_ ),
    .B1(\soc/simpleuart/_0382_ ),
    .Y(\soc/simpleuart/_0130_ ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1356_  (.CLK(clknet_leaf_92_clk),
    .D(net548),
    .Q(\soc/simpleuart_reg_div_do[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1357_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0001_ ),
    .Q(\soc/simpleuart_reg_div_do[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1358_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0002_ ),
    .Q(\soc/simpleuart_reg_div_do[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1359_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0003_ ),
    .Q(\soc/simpleuart_reg_div_do[27] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1360_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0004_ ),
    .Q(\soc/simpleuart_reg_div_do[28] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1361_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0005_ ),
    .Q(\soc/simpleuart_reg_div_do[29] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1362_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0006_ ),
    .Q(\soc/simpleuart_reg_div_do[30] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1363_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0007_ ),
    .Q(\soc/simpleuart_reg_div_do[31] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1364_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/simpleuart/_0008_ ),
    .Q(\soc/simpleuart_reg_div_do[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1365_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0009_ ),
    .Q(\soc/simpleuart_reg_div_do[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1366_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0010_ ),
    .Q(\soc/simpleuart_reg_div_do[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1367_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0011_ ),
    .Q(\soc/simpleuart_reg_div_do[19] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1368_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0012_ ),
    .Q(\soc/simpleuart_reg_div_do[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1369_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0013_ ),
    .Q(\soc/simpleuart_reg_div_do[21] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1370_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0014_ ),
    .Q(\soc/simpleuart_reg_div_do[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1371_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0015_ ),
    .Q(\soc/simpleuart_reg_div_do[23] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1372_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0016_ ),
    .Q(\soc/simpleuart_reg_div_do[8] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1373_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0017_ ),
    .Q(\soc/simpleuart_reg_div_do[9] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1374_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0018_ ),
    .Q(\soc/simpleuart_reg_div_do[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1375_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0019_ ),
    .Q(\soc/simpleuart_reg_div_do[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1376_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/simpleuart/_0020_ ),
    .Q(\soc/simpleuart_reg_div_do[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1377_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/simpleuart/_0021_ ),
    .Q(\soc/simpleuart_reg_div_do[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1378_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0022_ ),
    .Q(\soc/simpleuart_reg_div_do[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1379_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0023_ ),
    .Q(\soc/simpleuart_reg_div_do[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1380_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0024_ ),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1381_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0025_ ),
    .Q(\soc/simpleuart/send_pattern[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1382_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0026_ ),
    .Q(\soc/simpleuart/send_pattern[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1383_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0027_ ),
    .Q(\soc/simpleuart/send_pattern[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1384_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0028_ ),
    .Q(\soc/simpleuart/send_pattern[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1385_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0029_ ),
    .Q(\soc/simpleuart/send_pattern[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1386_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0030_ ),
    .Q(\soc/simpleuart/send_pattern[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1387_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0031_ ),
    .Q(\soc/simpleuart/send_pattern[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1388_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0032_ ),
    .Q(\soc/simpleuart/send_pattern[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1389_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0033_ ),
    .Q(\soc/simpleuart/send_bitcnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1390_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0034_ ),
    .Q(\soc/simpleuart/send_bitcnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1391_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0035_ ),
    .Q(\soc/simpleuart/send_bitcnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1392_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0036_ ),
    .Q(\soc/simpleuart/send_bitcnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1393_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0037_ ),
    .Q(\soc/simpleuart/send_dummy ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1394_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0038_ ),
    .Q(\soc/simpleuart/recv_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1395_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0039_ ),
    .Q(\soc/simpleuart/recv_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1396_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0040_ ),
    .Q(\soc/simpleuart/recv_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1397_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0041_ ),
    .Q(\soc/simpleuart/recv_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1398_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0042_ ),
    .Q(\soc/simpleuart/send_divcnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1399_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0043_ ),
    .Q(\soc/simpleuart/send_divcnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1400_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0044_ ),
    .Q(\soc/simpleuart/send_divcnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1401_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0045_ ),
    .Q(\soc/simpleuart/send_divcnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1402_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0046_ ),
    .Q(\soc/simpleuart/send_divcnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1403_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0047_ ),
    .Q(\soc/simpleuart/send_divcnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1404_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0048_ ),
    .Q(\soc/simpleuart/send_divcnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1405_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0049_ ),
    .Q(\soc/simpleuart/send_divcnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1406_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0050_ ),
    .Q(\soc/simpleuart/send_divcnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1407_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0051_ ),
    .Q(\soc/simpleuart/send_divcnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1408_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0052_ ),
    .Q(\soc/simpleuart/send_divcnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1409_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0053_ ),
    .Q(\soc/simpleuart/send_divcnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1410_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0054_ ),
    .Q(\soc/simpleuart/send_divcnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1411_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0055_ ),
    .Q(\soc/simpleuart/send_divcnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1412_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0056_ ),
    .Q(\soc/simpleuart/send_divcnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1413_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0057_ ),
    .Q(\soc/simpleuart/send_divcnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1414_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0058_ ),
    .Q(\soc/simpleuart/send_divcnt[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1415_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0059_ ),
    .Q(\soc/simpleuart/send_divcnt[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1416_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0060_ ),
    .Q(\soc/simpleuart/send_divcnt[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1417_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0061_ ),
    .Q(\soc/simpleuart/send_divcnt[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1418_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0062_ ),
    .Q(\soc/simpleuart/send_divcnt[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1419_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0063_ ),
    .Q(\soc/simpleuart/send_divcnt[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1420_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0064_ ),
    .Q(\soc/simpleuart/send_divcnt[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1421_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0065_ ),
    .Q(\soc/simpleuart/send_divcnt[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1422_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0066_ ),
    .Q(\soc/simpleuart/send_divcnt[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1423_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0067_ ),
    .Q(\soc/simpleuart/send_divcnt[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1424_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0068_ ),
    .Q(\soc/simpleuart/send_divcnt[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1425_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0069_ ),
    .Q(\soc/simpleuart/send_divcnt[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1426_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0070_ ),
    .Q(\soc/simpleuart/send_divcnt[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1427_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0071_ ),
    .Q(\soc/simpleuart/send_divcnt[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1428_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0072_ ),
    .Q(\soc/simpleuart/send_divcnt[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1429_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0073_ ),
    .Q(\soc/simpleuart/send_divcnt[31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1430_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0074_ ),
    .Q(\soc/simpleuart/recv_pattern[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1431_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0075_ ),
    .Q(\soc/simpleuart/recv_pattern[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1432_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0076_ ),
    .Q(\soc/simpleuart/recv_pattern[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1433_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0077_ ),
    .Q(\soc/simpleuart/recv_pattern[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1434_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0078_ ),
    .Q(\soc/simpleuart/recv_pattern[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1435_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0079_ ),
    .Q(\soc/simpleuart/recv_pattern[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1436_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0080_ ),
    .Q(\soc/simpleuart/recv_pattern[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1437_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0081_ ),
    .Q(\soc/simpleuart/recv_pattern[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1438_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0082_ ),
    .Q(\soc/simpleuart/recv_buf_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1439_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0083_ ),
    .Q(\soc/simpleuart/recv_buf_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1440_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0084_ ),
    .Q(\soc/simpleuart/recv_buf_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1441_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0085_ ),
    .Q(\soc/simpleuart/recv_buf_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1442_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0086_ ),
    .Q(\soc/simpleuart/recv_buf_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1443_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0087_ ),
    .Q(\soc/simpleuart/recv_buf_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1444_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0088_ ),
    .Q(\soc/simpleuart/recv_buf_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1445_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0089_ ),
    .Q(\soc/simpleuart/recv_buf_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1446_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0090_ ),
    .Q(\soc/simpleuart/recv_divcnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1447_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0091_ ),
    .Q(\soc/simpleuart/recv_divcnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1448_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0092_ ),
    .Q(\soc/simpleuart/recv_divcnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1449_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0093_ ),
    .Q(\soc/simpleuart/recv_divcnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1450_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0094_ ),
    .Q(\soc/simpleuart/recv_divcnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1451_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0095_ ),
    .Q(\soc/simpleuart/recv_divcnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1452_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0096_ ),
    .Q(\soc/simpleuart/recv_divcnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1453_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0097_ ),
    .Q(\soc/simpleuart/recv_divcnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1454_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0098_ ),
    .Q(\soc/simpleuart/recv_divcnt[8] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1455_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0099_ ),
    .Q(\soc/simpleuart/recv_divcnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1456_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0100_ ),
    .Q(\soc/simpleuart/recv_divcnt[10] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1457_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0101_ ),
    .Q(\soc/simpleuart/recv_divcnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1458_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0102_ ),
    .Q(\soc/simpleuart/recv_divcnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1459_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0103_ ),
    .Q(\soc/simpleuart/recv_divcnt[13] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1460_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0104_ ),
    .Q(\soc/simpleuart/recv_divcnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1461_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0105_ ),
    .Q(\soc/simpleuart/recv_divcnt[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1462_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0106_ ),
    .Q(\soc/simpleuart/recv_divcnt[16] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1463_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/simpleuart/_0107_ ),
    .Q(\soc/simpleuart/recv_divcnt[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1464_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/simpleuart/_0108_ ),
    .Q(\soc/simpleuart/recv_divcnt[18] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1465_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/simpleuart/_0109_ ),
    .Q(\soc/simpleuart/recv_divcnt[19] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1466_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0110_ ),
    .Q(\soc/simpleuart/recv_divcnt[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1467_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0111_ ),
    .Q(\soc/simpleuart/recv_divcnt[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1468_  (.CLK(clknet_leaf_92_clk),
    .D(net513),
    .Q(\soc/simpleuart/recv_divcnt[22] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1469_  (.CLK(clknet_leaf_92_clk),
    .D(net543),
    .Q(\soc/simpleuart/recv_divcnt[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1470_  (.CLK(clknet_leaf_92_clk),
    .D(net556),
    .Q(\soc/simpleuart/recv_divcnt[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1471_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0115_ ),
    .Q(\soc/simpleuart/recv_divcnt[25] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1472_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0116_ ),
    .Q(\soc/simpleuart/recv_divcnt[26] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1473_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/simpleuart/_0117_ ),
    .Q(\soc/simpleuart/recv_divcnt[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1474_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0118_ ),
    .Q(\soc/simpleuart/recv_divcnt[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1475_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0119_ ),
    .Q(\soc/simpleuart/recv_divcnt[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1476_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0120_ ),
    .Q(\soc/simpleuart/recv_divcnt[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1477_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/simpleuart/_0121_ ),
    .Q(\soc/simpleuart/recv_divcnt[31] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1478_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0122_ ),
    .Q(\soc/simpleuart_reg_div_do[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1479_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0123_ ),
    .Q(\soc/simpleuart_reg_div_do[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1480_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0124_ ),
    .Q(\soc/simpleuart_reg_div_do[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1481_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0125_ ),
    .Q(\soc/simpleuart_reg_div_do[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1482_  (.CLK(clknet_leaf_71_clk),
    .D(\soc/simpleuart/_0126_ ),
    .Q(\soc/simpleuart_reg_div_do[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1483_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0127_ ),
    .Q(\soc/simpleuart_reg_div_do[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/simpleuart/_1484_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0128_ ),
    .Q(\soc/simpleuart_reg_div_do[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/simpleuart/_1485_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/simpleuart/_0129_ ),
    .Q(\soc/simpleuart_reg_div_do[7] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/simpleuart/_1486_  (.CLK(clknet_leaf_76_clk),
    .D(\soc/simpleuart/_0130_ ),
    .Q(\soc/simpleuart/recv_buf_valid ));
 sky130_fd_sc_hd__xor2_2 \soc/spimemio/_0548_  (.A(\soc/spimemio/rd_addr[9] ),
    .B(net357),
    .X(\soc/spimemio/_0132_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0549_  (.A(\soc/spimemio/rd_addr[20] ),
    .B(\iomem_addr[20] ),
    .X(\soc/spimemio/_0133_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0550_  (.A(\soc/spimemio/rd_addr[21] ),
    .B(\iomem_addr[21] ),
    .X(\soc/spimemio/_0134_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0551_  (.A(\soc/spimemio/rd_addr[7] ),
    .B(net497),
    .X(\soc/spimemio/_0135_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0552_  (.A(\soc/spimemio/rd_addr[5] ),
    .B(net373),
    .X(\soc/spimemio/_0136_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0553_  (.A(net750),
    .B(net384),
    .X(\soc/spimemio/_0137_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0554_  (.A(\soc/spimemio/rd_addr[8] ),
    .B(net361),
    .Y(\soc/spimemio/_0138_ ));
 sky130_fd_sc_hd__nor4b_1 \soc/spimemio/_0555_  (.A(\soc/spimemio/_0135_ ),
    .B(\soc/spimemio/_0136_ ),
    .C(\soc/spimemio/_0137_ ),
    .D_N(\soc/spimemio/_0138_ ),
    .Y(\soc/spimemio/_0139_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0556_  (.A(net824),
    .B(\iomem_addr[13] ),
    .Y(\soc/spimemio/_0140_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0557_  (.A(\soc/spimemio/rd_addr[12] ),
    .B(net771),
    .Y(\soc/spimemio/_0141_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0559_  (.A(\soc/spimemio/rd_addr[15] ),
    .B(net713),
    .X(\soc/spimemio/_0143_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0560_  (.A(\soc/spimemio/rd_addr[19] ),
    .B(\iomem_addr[19] ),
    .X(\soc/spimemio/_0144_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0561_  (.A(\soc/spimemio/_0143_ ),
    .B(\soc/spimemio/_0144_ ),
    .Y(\soc/spimemio/_0145_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0562_  (.A(\soc/spimemio/_0139_ ),
    .B(net825),
    .C(\soc/spimemio/_0141_ ),
    .D(\soc/spimemio/_0145_ ),
    .Y(\soc/spimemio/_0146_ ));
 sky130_fd_sc_hd__or4_1 \soc/spimemio/_0563_  (.A(\soc/spimemio/_0132_ ),
    .B(\soc/spimemio/_0133_ ),
    .C(\soc/spimemio/_0134_ ),
    .D(net826),
    .X(\soc/spimemio/_0147_ ));
 sky130_fd_sc_hd__xnor2_2 \soc/spimemio/_0564_  (.A(\soc/spimemio/rd_addr[0] ),
    .B(net452),
    .Y(\soc/spimemio/_0148_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0565_  (.A(\soc/spimemio/rd_addr[1] ),
    .B(net453),
    .Y(\soc/spimemio/_0149_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0566_  (.A(\soc/spimemio/rd_addr[23] ),
    .Y(\soc/spimemio/_0150_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/spimemio/_0568_  (.A(net724),
    .SLEEP(net884),
    .X(\soc/spimemio/_0152_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/spimemio/_0569_  (.A(net392),
    .SLEEP(net747),
    .X(\soc/spimemio/_0153_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/spimemio/_0570_  (.A1(\soc/spimemio/_0150_ ),
    .A2(net694),
    .B1(\soc/spimemio/_0152_ ),
    .C1(\soc/spimemio/_0153_ ),
    .Y(\soc/spimemio/_0154_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0571_  (.A(\soc/spimemio/rd_addr[4] ),
    .Y(\soc/spimemio/_0155_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0572_  (.A(\soc/spimemio/rd_addr[14] ),
    .Y(\soc/spimemio/_0156_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0573_  (.A(net368),
    .Y(\soc/spimemio/_0157_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0574_  (.A(\soc/spimemio/rd_addr[10] ),
    .Y(\soc/spimemio/_0158_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0575_  (.A1(net783),
    .A2(\soc/spimemio/_0157_ ),
    .B1(\soc/spimemio/_0158_ ),
    .B2(net714),
    .Y(\soc/spimemio/_0159_ ));
 sky130_fd_sc_hd__a221oi_2 \soc/spimemio/_0576_  (.A1(\soc/spimemio/_0155_ ),
    .A2(net380),
    .B1(\soc/spimemio/_0156_ ),
    .B2(net708),
    .C1(\soc/spimemio/_0159_ ),
    .Y(\soc/spimemio/_0160_ ));
 sky130_fd_sc_hd__nand4_2 \soc/spimemio/_0577_  (.A(\soc/spimemio/_0148_ ),
    .B(\soc/spimemio/_0149_ ),
    .C(\soc/spimemio/_0154_ ),
    .D(\soc/spimemio/_0160_ ),
    .Y(\soc/spimemio/_0161_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0578_  (.A(net714),
    .Y(\soc/spimemio/_0162_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0579_  (.A(\soc/spimemio/rd_addr[17] ),
    .B(net779),
    .Y(\soc/spimemio/_0163_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/spimemio/_0580_  (.A1(\soc/spimemio/rd_addr[10] ),
    .A2(\soc/spimemio/_0162_ ),
    .B1(net822),
    .C1(\soc/spimemio/_0163_ ),
    .D1(net727),
    .Y(\soc/spimemio/_0164_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0581_  (.A(net728),
    .B(net736),
    .X(\soc/spimemio/_0165_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0582_  (.A(\soc/spimemio/rd_addr[11] ),
    .B(net744),
    .X(\soc/spimemio/_0166_ ));
 sky130_fd_sc_hd__or3_1 \soc/spimemio/_0583_  (.A(\soc/spimemio/_0164_ ),
    .B(\soc/spimemio/_0165_ ),
    .C(\soc/spimemio/_0166_ ),
    .X(\soc/spimemio/_0167_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0584_  (.A(net783),
    .Y(\soc/spimemio/_0168_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0585_  (.A1(\soc/spimemio/_0155_ ),
    .A2(net379),
    .B1(\soc/spimemio/_0168_ ),
    .B2(net369),
    .Y(\soc/spimemio/_0169_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0586_  (.A(\iomem_addr[22] ),
    .Y(\soc/spimemio/_0170_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \soc/spimemio/_0587_  (.A1_N(net864),
    .A2_N(\soc/spimemio/_0170_ ),
    .B1(\soc/spimemio/_0150_ ),
    .B2(net694),
    .Y(\soc/spimemio/_0171_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/spimemio/_0588_  (.A(net747),
    .SLEEP(net393),
    .X(\soc/spimemio/_0172_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/spimemio/_0589_  (.A(net884),
    .SLEEP(net724),
    .X(\soc/spimemio/_0173_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0590_  (.A(\soc/spimemio/_0172_ ),
    .B(\soc/spimemio/_0173_ ),
    .Y(\soc/spimemio/_0174_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/spimemio/_0591_  (.A1(\soc/spimemio/_0156_ ),
    .A2(net708),
    .B1(net864),
    .B2(\soc/spimemio/_0170_ ),
    .C1(\soc/spimemio/_0174_ ),
    .Y(\soc/spimemio/_0175_ ));
 sky130_fd_sc_hd__or4_1 \soc/spimemio/_0592_  (.A(\soc/spimemio/_0167_ ),
    .B(\soc/spimemio/_0169_ ),
    .C(\soc/spimemio/_0171_ ),
    .D(\soc/spimemio/_0175_ ),
    .X(\soc/spimemio/_0176_ ));
 sky130_fd_sc_hd__nor3_4 \soc/spimemio/_0593_  (.A(net827),
    .B(\soc/spimemio/_0161_ ),
    .C(\soc/spimemio/_0176_ ),
    .Y(\soc/spimem_ready ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0594_  (.A(\soc/spimemio/state[7] ),
    .Y(\soc/spimemio/_0177_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0595_  (.A(\soc/spimemio/rd_addr[9] ),
    .Y(\soc/spimemio/_0178_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0596_  (.A(\soc/spimemio/rd_addr[11] ),
    .Y(\soc/spimemio/_0179_ ));
 sky130_fd_sc_hd__and4_2 \soc/spimemio/_0597_  (.A(net747),
    .B(net750),
    .C(\soc/spimemio/rd_addr[4] ),
    .D(\soc/spimemio/rd_addr[5] ),
    .X(\soc/spimemio/_0180_ ));
 sky130_fd_sc_hd__nand4_2 \soc/spimemio/_0598_  (.A(\soc/spimemio/rd_addr[6] ),
    .B(\soc/spimemio/rd_addr[7] ),
    .C(\soc/spimemio/rd_addr[8] ),
    .D(\soc/spimemio/_0180_ ),
    .Y(\soc/spimemio/_0181_ ));
 sky130_fd_sc_hd__nor4_2 \soc/spimemio/_0599_  (.A(\soc/spimemio/_0178_ ),
    .B(\soc/spimemio/_0158_ ),
    .C(\soc/spimemio/_0179_ ),
    .D(\soc/spimemio/_0181_ ),
    .Y(\soc/spimemio/_0182_ ));
 sky130_fd_sc_hd__and4_4 \soc/spimemio/_0600_  (.A(\soc/spimemio/rd_addr[12] ),
    .B(\soc/spimemio/rd_addr[13] ),
    .C(\soc/spimemio/rd_addr[14] ),
    .D(\soc/spimemio/_0182_ ),
    .X(\soc/spimemio/_0183_ ));
 sky130_fd_sc_hd__and4_2 \soc/spimemio/_0601_  (.A(\soc/spimemio/rd_addr[15] ),
    .B(net728),
    .C(\soc/spimemio/rd_addr[17] ),
    .D(\soc/spimemio/_0183_ ),
    .X(\soc/spimemio/_0184_ ));
 sky130_fd_sc_hd__and4_2 \soc/spimemio/_0603_  (.A(\soc/spimemio/rd_addr[18] ),
    .B(\soc/spimemio/rd_addr[19] ),
    .C(\soc/spimemio/rd_addr[20] ),
    .D(\soc/spimemio/_0184_ ),
    .X(\soc/spimemio/_0186_ ));
 sky130_fd_sc_hd__and2_1 \soc/spimemio/_0605_  (.A(\soc/spimemio/rd_addr[21] ),
    .B(\soc/spimemio/_0186_ ),
    .X(\soc/spimemio/_0188_ ));
 sky130_fd_sc_hd__xnor3_1 \soc/spimemio/_0606_  (.A(\soc/spimemio/rd_addr[22] ),
    .B(\soc/spimemio/_0170_ ),
    .C(\soc/spimemio/_0188_ ),
    .X(\soc/spimemio/_0189_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_0607_  (.A1(net939),
    .A2(net864),
    .A3(\soc/spimemio/_0186_ ),
    .B1(\soc/spimemio/rd_addr[23] ),
    .Y(\soc/spimemio/_0190_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0608_  (.A(net694),
    .B(\soc/spimemio/_0190_ ),
    .Y(\soc/spimemio/_0191_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0609_  (.A(net939),
    .B(net864),
    .C(\soc/spimemio/rd_addr[23] ),
    .D(\soc/spimemio/_0186_ ),
    .Y(\soc/spimemio/_0192_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0610_  (.A(\soc/spimemio/_0134_ ),
    .B(\soc/spimemio/_0186_ ),
    .Y(\soc/spimemio/_0193_ ));
 sky130_fd_sc_hd__a41oi_1 \soc/spimemio/_0612_  (.A1(\soc/spimemio/rd_addr[15] ),
    .A2(net728),
    .A3(\soc/spimemio/rd_addr[17] ),
    .A4(\soc/spimemio/_0183_ ),
    .B1(\soc/spimemio/_0173_ ),
    .Y(\soc/spimemio/_0195_ ));
 sky130_fd_sc_hd__o21bai_1 \soc/spimemio/_0613_  (.A1(\soc/spimemio/_0152_ ),
    .A2(\soc/spimemio/_0195_ ),
    .B1_N(\soc/spimemio/_0144_ ),
    .Y(\soc/spimemio/_0196_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0614_  (.A(\soc/spimemio/rd_addr[18] ),
    .B(\soc/spimemio/_0144_ ),
    .C(\soc/spimemio/_0184_ ),
    .Y(\soc/spimemio/_0197_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0615_  (.A(\soc/spimemio/rd_addr[18] ),
    .B(\soc/spimemio/_0184_ ),
    .Y(\soc/spimemio/_0198_ ));
 sky130_fd_sc_hd__a22oi_2 \soc/spimemio/_0616_  (.A1(\soc/spimemio/_0196_ ),
    .A2(\soc/spimemio/_0197_ ),
    .B1(\soc/spimemio/_0198_ ),
    .B2(net724),
    .Y(\soc/spimemio/_0199_ ));
 sky130_fd_sc_hd__a31o_1 \soc/spimemio/_0617_  (.A1(\soc/spimemio/rd_addr[18] ),
    .A2(\soc/spimemio/rd_addr[19] ),
    .A3(\soc/spimemio/_0184_ ),
    .B1(\soc/spimemio/_0133_ ),
    .X(\soc/spimemio/_0200_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0618_  (.A(\soc/spimemio/rd_addr[18] ),
    .B(\soc/spimemio/rd_addr[19] ),
    .C(\soc/spimemio/_0133_ ),
    .D(\soc/spimemio/_0184_ ),
    .Y(\soc/spimemio/_0201_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0619_  (.A(\soc/spimemio/rd_addr[15] ),
    .B(net728),
    .C(\soc/spimemio/_0183_ ),
    .X(\soc/spimemio/_0202_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0620_  (.A(\soc/spimemio/_0163_ ),
    .B(\soc/spimemio/_0202_ ),
    .Y(\soc/spimemio/_0203_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0621_  (.A1(\soc/spimemio/rd_addr[15] ),
    .A2(\soc/spimemio/_0183_ ),
    .B1(\soc/spimemio/_0165_ ),
    .Y(\soc/spimemio/_0204_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0622_  (.A(\soc/spimemio/rd_addr[15] ),
    .B(\soc/spimemio/_0165_ ),
    .C(\soc/spimemio/_0183_ ),
    .X(\soc/spimemio/_0205_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0623_  (.A(\soc/spimemio/rd_addr[12] ),
    .B(\soc/spimemio/rd_addr[13] ),
    .C(\soc/spimemio/_0182_ ),
    .X(\soc/spimemio/_0206_ ));
 sky130_fd_sc_hd__xnor3_1 \soc/spimemio/_0624_  (.A(\soc/spimemio/rd_addr[14] ),
    .B(net708),
    .C(\soc/spimemio/_0206_ ),
    .X(\soc/spimemio/_0207_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/spimemio/_0625_  (.A1(\soc/spimemio/_0204_ ),
    .A2(\soc/spimemio/_0205_ ),
    .B1(\soc/spimemio/_0207_ ),
    .Y(\soc/spimemio/_0208_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0626_  (.A(\soc/spimemio/_0143_ ),
    .B(\soc/spimemio/_0183_ ),
    .Y(\soc/spimemio/_0209_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0627_  (.A(\soc/spimemio/rd_addr[15] ),
    .B(net728),
    .C(\soc/spimemio/_0163_ ),
    .D(\soc/spimemio/_0183_ ),
    .Y(\soc/spimemio/_0210_ ));
 sky130_fd_sc_hd__and4_1 \soc/spimemio/_0628_  (.A(\soc/spimemio/rd_addr[6] ),
    .B(\soc/spimemio/rd_addr[7] ),
    .C(\soc/spimemio/rd_addr[8] ),
    .D(\soc/spimemio/_0180_ ),
    .X(\soc/spimemio/_0211_ ));
 sky130_fd_sc_hd__nand3_2 \soc/spimemio/_0629_  (.A(\soc/spimemio/rd_addr[9] ),
    .B(\soc/spimemio/rd_addr[10] ),
    .C(\soc/spimemio/_0211_ ),
    .Y(\soc/spimemio/_0212_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0630_  (.A(\soc/spimemio/_0166_ ),
    .B(\soc/spimemio/_0212_ ),
    .Y(\soc/spimemio/_0213_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0631_  (.A(\soc/spimemio/rd_addr[6] ),
    .B(\soc/spimemio/_0180_ ),
    .Y(\soc/spimemio/_0214_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0632_  (.A(\soc/spimemio/_0157_ ),
    .B(\soc/spimemio/_0214_ ),
    .Y(\soc/spimemio/_0215_ ));
 sky130_fd_sc_hd__and2_1 \soc/spimemio/_0633_  (.A(\soc/spimemio/rd_addr[6] ),
    .B(\soc/spimemio/_0180_ ),
    .X(\soc/spimemio/_0216_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0634_  (.A(\soc/spimemio/_0135_ ),
    .B(\soc/spimemio/_0216_ ),
    .Y(\soc/spimemio/_0217_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0635_  (.A(net747),
    .B(\soc/spimemio/rd_addr[3] ),
    .C(\soc/spimemio/rd_addr[4] ),
    .Y(\soc/spimemio/_0218_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0636_  (.A(\soc/spimemio/_0136_ ),
    .B(\soc/spimemio/_0218_ ),
    .X(\soc/spimemio/_0219_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0637_  (.A(\soc/spimemio/_0148_ ),
    .B(\soc/spimemio/_0149_ ),
    .C(\soc/spimemio/_0219_ ),
    .X(\soc/spimemio/_0220_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0638_  (.A(\soc/spimemio/_0215_ ),
    .B(\soc/spimemio/_0217_ ),
    .C(\soc/spimemio/_0220_ ),
    .Y(\soc/spimemio/_0221_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0639_  (.A(\soc/spimemio/rd_addr[6] ),
    .B(\soc/spimemio/rd_addr[7] ),
    .C(\soc/spimemio/_0180_ ),
    .X(\soc/spimemio/_0222_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0640_  (.A(net747),
    .B(net750),
    .Y(\soc/spimemio/_0223_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0641_  (.A(\soc/spimemio/_0155_ ),
    .B(\soc/spimemio/_0223_ ),
    .Y(\soc/spimemio/_0224_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/_0642_  (.A(net377),
    .B(\soc/spimemio/_0224_ ),
    .X(\soc/spimemio/_0225_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0643_  (.A(\soc/spimemio/_0132_ ),
    .B(\soc/spimemio/_0211_ ),
    .Y(\soc/spimemio/_0226_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/spimemio/_0644_  (.A0(\soc/spimemio/_0153_ ),
    .A1(\soc/spimemio/_0172_ ),
    .S(\soc/spimemio/_0137_ ),
    .Y(\soc/spimemio/_0227_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0645_  (.A1(\soc/spimemio/_0138_ ),
    .A2(\soc/spimemio/_0222_ ),
    .B1(\soc/spimemio/_0227_ ),
    .Y(\soc/spimemio/_0228_ ));
 sky130_fd_sc_hd__o2111ai_1 \soc/spimemio/_0646_  (.A1(\soc/spimemio/_0138_ ),
    .A2(\soc/spimemio/_0222_ ),
    .B1(\soc/spimemio/_0225_ ),
    .C1(\soc/spimemio/_0226_ ),
    .D1(\soc/spimemio/_0228_ ),
    .Y(\soc/spimemio/_0229_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0647_  (.A(\soc/spimemio/_0213_ ),
    .B(\soc/spimemio/_0221_ ),
    .C(\soc/spimemio/_0229_ ),
    .Y(\soc/spimemio/_0230_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/spimemio/_0648_  (.A1(\soc/spimemio/_0178_ ),
    .A2(\soc/spimemio/_0181_ ),
    .B1(\soc/spimemio/_0158_ ),
    .Y(\soc/spimemio/_0231_ ));
 sky130_fd_sc_hd__a21o_1 \soc/spimemio/_0649_  (.A1(\soc/spimemio/_0212_ ),
    .A2(\soc/spimemio/_0231_ ),
    .B1(net714),
    .X(\soc/spimemio/_0232_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0650_  (.A(net714),
    .B(\soc/spimemio/_0212_ ),
    .C(\soc/spimemio/_0231_ ),
    .Y(\soc/spimemio/_0233_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0651_  (.A(\soc/spimemio/_0141_ ),
    .B(\soc/spimemio/_0182_ ),
    .Y(\soc/spimemio/_0234_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0652_  (.A1(\soc/spimemio/rd_addr[12] ),
    .A2(\soc/spimemio/_0182_ ),
    .B1(\soc/spimemio/_0140_ ),
    .Y(\soc/spimemio/_0235_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0653_  (.A(\soc/spimemio/rd_addr[12] ),
    .B(\soc/spimemio/_0140_ ),
    .C(\soc/spimemio/_0182_ ),
    .X(\soc/spimemio/_0236_ ));
 sky130_fd_sc_hd__a2111oi_1 \soc/spimemio/_0654_  (.A1(\soc/spimemio/_0232_ ),
    .A2(\soc/spimemio/_0233_ ),
    .B1(\soc/spimemio/_0234_ ),
    .C1(\soc/spimemio/_0235_ ),
    .D1(\soc/spimemio/_0236_ ),
    .Y(\soc/spimemio/_0237_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0655_  (.A(\soc/spimemio/_0209_ ),
    .B(net729),
    .C(\soc/spimemio/_0230_ ),
    .D(\soc/spimemio/_0237_ ),
    .Y(\soc/spimemio/_0238_ ));
 sky130_fd_sc_hd__a2111oi_1 \soc/spimemio/_0656_  (.A1(\soc/spimemio/_0200_ ),
    .A2(\soc/spimemio/_0201_ ),
    .B1(\soc/spimemio/_0203_ ),
    .C1(\soc/spimemio/_0208_ ),
    .D1(net730),
    .Y(\soc/spimemio/_0239_ ));
 sky130_fd_sc_hd__nand4_2 \soc/spimemio/_0657_  (.A(\soc/spimemio/_0192_ ),
    .B(\soc/spimemio/_0193_ ),
    .C(\soc/spimemio/_0199_ ),
    .D(net731),
    .Y(\soc/spimemio/_0240_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0658_  (.A(net822),
    .Y(\soc/spimemio/_0241_ ));
 sky130_fd_sc_hd__nand2b_2 \soc/spimemio/_0659_  (.A_N(\soc/spimem_ready ),
    .B(net727),
    .Y(\soc/spimemio/_0242_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0660_  (.A(\soc/spimemio/_0241_ ),
    .B(\soc/spimemio/_0242_ ),
    .Y(\soc/spimemio/_0243_ ));
 sky130_fd_sc_hd__o31ai_4 \soc/spimemio/_0661_  (.A1(net865),
    .A2(\soc/spimemio/_0191_ ),
    .A3(net732),
    .B1(\soc/spimemio/_0243_ ),
    .Y(\soc/spimemio/_0244_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_8 \soc/spimemio/_0662_  (.A(_074_),
    .SLEEP(net735),
    .X(\soc/spimemio/_0245_ ));
 sky130_fd_sc_hd__nand2_2 \soc/spimemio/_0663_  (.A(net733),
    .B(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0246_ ));
 sky130_fd_sc_hd__nand3_4 \soc/spimemio/_0665_  (.A(\soc/spimemio/xfer/_047_ ),
    .B(net733),
    .C(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0248_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0666_  (.A(\soc/spimemio/state[0] ),
    .Y(\soc/spimemio/_0249_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/spimemio/_0667_  (.A1(\soc/spimemio/dout_valid ),
    .A2(\soc/spimemio/_0177_ ),
    .A3(\soc/spimemio/_0246_ ),
    .B1(\soc/spimemio/_0248_ ),
    .B2(\soc/spimemio/_0249_ ),
    .Y(\soc/spimemio/_0010_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/spimemio/_0669_  (.A(\soc/spimemio/state[9] ),
    .SLEEP(\soc/spimemio/_0242_ ),
    .X(\soc/spimemio/_0251_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0670_  (.A(\soc/spimemio/_0251_ ),
    .Y(\soc/spimemio/_0252_ ));
 sky130_fd_sc_hd__nand2b_4 \soc/spimemio/_0673_  (.A_N(\soc/spimemio/softreset ),
    .B(_074_),
    .Y(\soc/spimemio/_0255_ ));
 sky130_fd_sc_hd__nor2_2 \soc/spimemio/_0675_  (.A(\soc/spimemio/xfer/_047_ ),
    .B(\soc/spimemio/_0255_ ),
    .Y(\soc/spimemio/_0257_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0676_  (.A(\soc/spimemio/state[6] ),
    .B(net733),
    .C(\soc/spimemio/_0257_ ),
    .Y(\soc/spimemio/_0258_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0677_  (.A1(\soc/spimemio/_0248_ ),
    .A2(\soc/spimemio/_0252_ ),
    .B1(\soc/spimemio/_0258_ ),
    .Y(\soc/spimemio/_0009_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0678_  (.A(\soc/spimemio/state[8] ),
    .Y(\soc/spimemio/_0259_ ));
 sky130_fd_sc_hd__nand2_2 \soc/spimemio/_0679_  (.A(net733),
    .B(\soc/spimemio/_0257_ ),
    .Y(\soc/spimemio/_0260_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0680_  (.A(\soc/spimemio/state[5] ),
    .Y(\soc/spimemio/_0261_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0681_  (.A1(\soc/spimemio/_0259_ ),
    .A2(\soc/spimemio/_0248_ ),
    .B1(\soc/spimemio/_0260_ ),
    .B2(\soc/spimemio/_0261_ ),
    .Y(\soc/spimemio/_0008_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0682_  (.A(\soc/spimemio/dout_valid ),
    .Y(\soc/spimemio/_0262_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0683_  (.A(\soc/spimemio/state[4] ),
    .Y(\soc/spimemio/_0263_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/spimemio/_0684_  (.A1(\soc/spimemio/_0262_ ),
    .A2(\soc/spimemio/_0177_ ),
    .A3(\soc/spimemio/_0246_ ),
    .B1(\soc/spimemio/_0260_ ),
    .B2(\soc/spimemio/_0263_ ),
    .Y(\soc/spimemio/_0007_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0685_  (.A(\soc/spimemio/state[11] ),
    .Y(\soc/spimemio/_0264_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/spimemio/_0686_  (.A_N(net727),
    .B(\soc/spimemio/rd_wait ),
    .C(\soc/spimemio/state[3] ),
    .Y(\soc/spimemio/_0265_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/_0687_  (.A_N(net727),
    .B(\soc/spimemio/rd_wait ),
    .Y(\soc/spimemio/_0266_ ));
 sky130_fd_sc_hd__and2_0 \soc/spimemio/_0688_  (.A(\soc/spimemio/state[3] ),
    .B(\soc/spimemio/_0266_ ),
    .X(\soc/spimemio/_0267_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0689_  (.A(net733),
    .B(\soc/spimemio/_0257_ ),
    .C(\soc/spimemio/_0267_ ),
    .Y(\soc/spimemio/_0268_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/spimemio/_0690_  (.A1(\soc/spimemio/_0264_ ),
    .A2(\soc/spimemio/_0248_ ),
    .B1(\soc/spimemio/_0265_ ),
    .B2(\soc/spimemio/_0246_ ),
    .C1(\soc/spimemio/_0268_ ),
    .Y(\soc/spimemio/_0006_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0691_  (.A(\soc/spimemio/state[2] ),
    .Y(\soc/spimemio/_0269_ ));
 sky130_fd_sc_hd__or2_0 \soc/spimemio/_0692_  (.A(net746),
    .B(net733),
    .X(\soc/spimemio/_0270_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0694_  (.A(\soc/spimemio/dout_valid ),
    .B(\soc/spimemio/state[10] ),
    .C(net733),
    .D(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0272_ ));
 sky130_fd_sc_hd__o221ai_1 \soc/spimemio/_0695_  (.A1(\soc/spimemio/_0269_ ),
    .A2(\soc/spimemio/_0260_ ),
    .B1(\soc/spimemio/_0270_ ),
    .B2(\soc/spimemio/_0255_ ),
    .C1(\soc/spimemio/_0272_ ),
    .Y(\soc/spimemio/_0005_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0696_  (.A(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/_0273_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0697_  (.A(\soc/spimemio/_0273_ ),
    .B(\soc/spimemio/state[1] ),
    .Y(\soc/spimemio/_0274_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0699_  (.A1(\soc/spimemio/config_ddr ),
    .A2(\soc/spimemio/config_qspi ),
    .B1(\soc/spimemio/state[12] ),
    .Y(\soc/spimemio/_0276_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0700_  (.A1(\soc/spimemio/_0246_ ),
    .A2(\soc/spimemio/_0274_ ),
    .B1(\soc/spimemio/_0276_ ),
    .B2(\soc/spimemio/_0248_ ),
    .Y(\soc/spimemio/_0004_ ));
 sky130_fd_sc_hd__a31o_1 \soc/spimemio/_0701_  (.A1(\soc/spimemio/_0273_ ),
    .A2(\soc/spimemio/state[0] ),
    .A3(net733),
    .B1(\soc/spimemio/_0255_ ),
    .X(\soc/spimemio/_0000_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \soc/spimemio/_0702_  (.A(\soc/spimemio/state[12] ),
    .SLEEP(\soc/spimemio/xfer/_047_ ),
    .X(\soc/spimemio/_0277_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0703_  (.A1(\soc/spimemio/xfer/_047_ ),
    .A2(\soc/spimemio/state[6] ),
    .B1(\soc/spimemio/_0277_ ),
    .Y(\soc/spimemio/_0278_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0704_  (.A(\soc/spimemio/_0246_ ),
    .B(\soc/spimemio/_0278_ ),
    .Y(\soc/spimemio/_0003_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0705_  (.A1(\soc/spimemio/_0261_ ),
    .A2(\soc/spimemio/_0248_ ),
    .B1(\soc/spimemio/_0260_ ),
    .B2(\soc/spimemio/_0264_ ),
    .Y(\soc/spimemio/_0002_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0706_  (.A(\soc/spimemio/config_cont ),
    .Y(\soc/spimemio/_0279_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0707_  (.A(\soc/spimemio/state[9] ),
    .B(\soc/spimemio/_0242_ ),
    .Y(\soc/spimemio/_0280_ ));
 sky130_fd_sc_hd__o21a_1 \soc/spimemio/_0708_  (.A1(\soc/spimemio/_0279_ ),
    .A2(net733),
    .B1(\soc/spimemio/_0280_ ),
    .X(\soc/spimemio/_0281_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0709_  (.A(\soc/spimemio/xfer/_047_ ),
    .B(\soc/spimemio/state[2] ),
    .C(\soc/spimemio/_0244_ ),
    .D(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0282_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0710_  (.A(net733),
    .B(\soc/spimemio/_0257_ ),
    .C(\soc/spimemio/_0251_ ),
    .Y(\soc/spimemio/_0283_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/spimemio/_0711_  (.A1(\soc/spimemio/_0255_ ),
    .A2(\soc/spimemio/_0281_ ),
    .B1(\soc/spimemio/_0282_ ),
    .C1(\soc/spimemio/_0283_ ),
    .Y(\soc/spimemio/_0012_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0712_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/config_qspi ),
    .Y(\soc/spimemio/_0284_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/spimemio/_0713_  (.A1(\soc/spimemio/state[12] ),
    .A2(\soc/spimemio/_0284_ ),
    .B1(\soc/spimemio/_0267_ ),
    .C1(\soc/spimemio/state[1] ),
    .Y(\soc/spimemio/_0285_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0714_  (.A1(\soc/spimemio/_0259_ ),
    .A2(\soc/spimemio/_0260_ ),
    .B1(\soc/spimemio/_0285_ ),
    .B2(\soc/spimemio/_0248_ ),
    .Y(\soc/spimemio/_0011_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0715_  (.A(\soc/spimemio/_0262_ ),
    .B(\soc/spimemio/state[10] ),
    .C(net733),
    .D(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0286_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0716_  (.A1(\soc/spimemio/_0263_ ),
    .A2(\soc/spimemio/_0248_ ),
    .B1(\soc/spimemio/_0286_ ),
    .Y(\soc/spimemio/_0001_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \soc/spimemio/_0717_  (.A(\soc/spimemio/din_ddr ),
    .SLEEP(\soc/spimemio/din_qspi ),
    .X(\soc/spimemio/xfer_dspi ));
 sky130_fd_sc_hd__and2_0 \soc/spimemio/_0718_  (.A(\soc/spimemio/din_ddr ),
    .B(\soc/spimemio/din_qspi ),
    .X(\soc/spimemio/xfer_ddr ));
 sky130_fd_sc_hd__mux2_4 \soc/spimemio/_0721_  (.A0(\soc/spimemio/config_csb ),
    .A1(\soc/spimemio/xfer_csb ),
    .S(\soc/spimemio/config_en ),
    .X(net3));
 sky130_fd_sc_hd__mux2_4 \soc/spimemio/_0722_  (.A0(\soc/spimemio/config_clk ),
    .A1(\soc/spimemio/xfer_clk ),
    .S(\soc/spimemio/config_en ),
    .X(net2));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0723_  (.A0(\soc/spimemio/config_oe[0] ),
    .A1(\soc/spimemio/xfer_io0_oe ),
    .S(\soc/spimemio/config_en ),
    .X(flash_io0_oe));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0724_  (.A0(\soc/spimemio/config_oe[1] ),
    .A1(\soc/spimemio/xfer_io1_oe ),
    .S(\soc/spimemio/config_en ),
    .X(flash_io1_oe));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0725_  (.A0(\soc/spimemio/config_oe[2] ),
    .A1(\soc/spimemio/xfer_io2_oe ),
    .S(\soc/spimemio/config_en ),
    .X(flash_io2_oe));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0726_  (.A0(\soc/spimemio/config_oe[3] ),
    .A1(\soc/spimemio/xfer_io2_oe ),
    .S(\soc/spimemio/config_en ),
    .X(flash_io3_oe));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/_0727_  (.A_N(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io0_do ),
    .Y(\soc/spimemio/_0289_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0728_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io0_90 ),
    .Y(\soc/spimemio/_0290_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0729_  (.A(\soc/spimemio/config_en ),
    .B(\soc/spimemio/config_do[0] ),
    .Y(\soc/spimemio/_0291_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/spimemio/_0730_  (.A1(\soc/spimemio/config_en ),
    .A2(\soc/spimemio/_0289_ ),
    .A3(\soc/spimemio/_0290_ ),
    .B1(\soc/spimemio/_0291_ ),
    .Y(flash_io0));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/_0731_  (.A_N(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io1_do ),
    .Y(\soc/spimemio/_0292_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0732_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io1_90 ),
    .Y(\soc/spimemio/_0293_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0733_  (.A(\soc/spimemio/config_en ),
    .B(\soc/spimemio/config_do[1] ),
    .Y(\soc/spimemio/_0294_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/spimemio/_0734_  (.A1(\soc/spimemio/config_en ),
    .A2(\soc/spimemio/_0292_ ),
    .A3(\soc/spimemio/_0293_ ),
    .B1(\soc/spimemio/_0294_ ),
    .Y(flash_io1));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/_0735_  (.A_N(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io2_do ),
    .Y(\soc/spimemio/_0295_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0736_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io2_90 ),
    .Y(\soc/spimemio/_0296_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0737_  (.A(\soc/spimemio/config_en ),
    .B(\soc/spimemio/config_do[2] ),
    .Y(\soc/spimemio/_0297_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/spimemio/_0738_  (.A1(\soc/spimemio/config_en ),
    .A2(\soc/spimemio/_0295_ ),
    .A3(\soc/spimemio/_0296_ ),
    .B1(\soc/spimemio/_0297_ ),
    .Y(flash_io2));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/_0739_  (.A_N(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io3_do ),
    .Y(\soc/spimemio/_0298_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0740_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/xfer_io3_90 ),
    .Y(\soc/spimemio/_0299_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0741_  (.A(\soc/spimemio/config_en ),
    .B(\soc/spimemio/config_do[3] ),
    .Y(\soc/spimemio/_0300_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/spimemio/_0742_  (.A1(\soc/spimemio/config_en ),
    .A2(\soc/spimemio/_0298_ ),
    .A3(\soc/spimemio/_0299_ ),
    .B1(\soc/spimemio/_0300_ ),
    .Y(flash_io3));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0744_  (.A(\soc/spimemio/dout_tag[1] ),
    .B(\soc/spimemio/dout_tag[0] ),
    .C(\soc/spimemio/dout_valid ),
    .Y(\soc/spimemio/_0301_ ));
 sky130_fd_sc_hd__nor4_4 \soc/spimemio/_0745_  (.A(\soc/spimemio/dout_tag[3] ),
    .B(net722),
    .C(\soc/spimemio/_0255_ ),
    .D(\soc/spimemio/_0301_ ),
    .Y(\soc/spimemio/_0302_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0746_  (.A0(\soc/spimemio/buffer[16] ),
    .A1(\soc/spimemio/dout_data[0] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0014_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0747_  (.A0(\soc/spimemio/buffer[17] ),
    .A1(net753),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0015_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0748_  (.A0(\soc/spimemio/buffer[18] ),
    .A1(\soc/spimemio/dout_data[2] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0016_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0749_  (.A0(\soc/spimemio/buffer[19] ),
    .A1(\soc/spimemio/dout_data[3] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0017_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0750_  (.A0(\soc/spimemio/buffer[20] ),
    .A1(\soc/spimemio/dout_data[4] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0018_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0751_  (.A0(\soc/spimemio/buffer[21] ),
    .A1(\soc/spimemio/dout_data[5] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0019_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0752_  (.A0(\soc/spimemio/buffer[22] ),
    .A1(\soc/spimemio/dout_data[6] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0020_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0753_  (.A0(\soc/spimemio/buffer[23] ),
    .A1(\soc/spimemio/dout_data[7] ),
    .S(\soc/spimemio/_0302_ ),
    .X(\soc/spimemio/_0021_ ));
 sky130_fd_sc_hd__nor2_2 \soc/spimemio/_0754_  (.A(\soc/spimemio/dout_tag[0] ),
    .B(\soc/spimemio/_0262_ ),
    .Y(\soc/spimemio/_0303_ ));
 sky130_fd_sc_hd__nor2_2 \soc/spimemio/_0755_  (.A(\soc/spimemio/dout_tag[1] ),
    .B(\soc/spimemio/dout_tag[3] ),
    .Y(\soc/spimemio/_0304_ ));
 sky130_fd_sc_hd__nand4_4 \soc/spimemio/_0756_  (.A(net722),
    .B(\soc/spimemio/_0245_ ),
    .C(\soc/spimemio/_0303_ ),
    .D(\soc/spimemio/_0304_ ),
    .Y(\soc/spimemio/_0305_ ));
 sky130_fd_sc_hd__nor2_8 \soc/spimemio/_0757_  (.A(\soc/spimemio/rd_inc ),
    .B(net106),
    .Y(\soc/spimemio/_0306_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0759_  (.A(net454),
    .B(\soc/spimemio/_0306_ ),
    .Y(\soc/spimemio/_0308_ ));
 sky130_fd_sc_hd__or2_4 \soc/spimemio/_0760_  (.A(\soc/spimemio/rd_inc ),
    .B(net106),
    .X(\soc/spimemio/_0309_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0762_  (.A(\soc/spimemio/rd_addr[0] ),
    .B(\soc/spimemio/_0309_ ),
    .Y(\soc/spimemio/_0311_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0763_  (.A(\soc/spimemio/_0308_ ),
    .B(\soc/spimemio/_0311_ ),
    .Y(\soc/spimemio/_0025_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0764_  (.A(net455),
    .B(\soc/spimemio/_0306_ ),
    .Y(\soc/spimemio/_0312_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0765_  (.A(\soc/spimemio/rd_addr[1] ),
    .B(\soc/spimemio/_0309_ ),
    .Y(\soc/spimemio/_0313_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0766_  (.A(\soc/spimemio/_0312_ ),
    .B(\soc/spimemio/_0313_ ),
    .Y(\soc/spimemio/_0026_ ));
 sky130_fd_sc_hd__nand3_4 \soc/spimemio/_0768_  (.A(net722),
    .B(\soc/spimemio/_0303_ ),
    .C(\soc/spimemio/_0304_ ),
    .Y(\soc/spimemio/_0315_ ));
 sky130_fd_sc_hd__nor2_8 \soc/spimemio/_0769_  (.A(\soc/spimemio/_0255_ ),
    .B(\soc/spimemio/_0315_ ),
    .Y(\soc/spimemio/_0316_ ));
 sky130_fd_sc_hd__nand2_8 \soc/spimemio/_0770_  (.A(\soc/spimemio/rd_inc ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0317_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0772_  (.A(\soc/spimemio/rd_addr[2] ),
    .B(\soc/spimemio/_0317_ ),
    .Y(\soc/spimemio/_0319_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0773_  (.A1(\soc/spimemio/rd_addr[2] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(net390),
    .C1(\soc/spimemio/_0319_ ),
    .X(\soc/spimemio/_0027_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0774_  (.A(\soc/spimemio/rd_addr[2] ),
    .B(\soc/spimemio/rd_addr[3] ),
    .Y(\soc/spimemio/_0320_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \soc/spimemio/_0775_  (.A(\soc/spimemio/rd_inc ),
    .SLEEP(net106),
    .X(\soc/spimemio/_0321_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0776_  (.A1(\soc/spimemio/rd_addr[3] ),
    .A2(net106),
    .B1(\soc/spimemio/_0321_ ),
    .B2(\soc/spimemio/_0223_ ),
    .Y(\soc/spimemio/_0322_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0777_  (.A(net383),
    .B(\soc/spimemio/_0306_ ),
    .Y(\soc/spimemio/_0323_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0778_  (.A1(\soc/spimemio/_0320_ ),
    .A2(\soc/spimemio/_0322_ ),
    .B1(\soc/spimemio/_0323_ ),
    .Y(\soc/spimemio/_0028_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0780_  (.A(net376),
    .B(\soc/spimemio/_0309_ ),
    .Y(\soc/spimemio/_0325_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/spimemio/_0781_  (.A1(\soc/spimemio/_0155_ ),
    .A2(net106),
    .B1(\soc/spimemio/_0321_ ),
    .B2(\soc/spimemio/_0224_ ),
    .C1(\soc/spimemio/_0325_ ),
    .Y(\soc/spimemio/_0029_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0782_  (.A(net372),
    .B(\soc/spimemio/_0309_ ),
    .Y(\soc/spimemio/_0326_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0783_  (.A1(\soc/spimemio/rd_inc ),
    .A2(net748),
    .B1(net106),
    .Y(\soc/spimemio/_0327_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0784_  (.A(\soc/spimemio/rd_addr[5] ),
    .B(\soc/spimemio/_0327_ ),
    .Y(\soc/spimemio/_0328_ ));
 sky130_fd_sc_hd__a211oi_1 \soc/spimemio/_0785_  (.A1(\soc/spimemio/_0180_ ),
    .A2(\soc/spimemio/_0321_ ),
    .B1(\soc/spimemio/_0326_ ),
    .C1(\soc/spimemio/_0328_ ),
    .Y(\soc/spimemio/_0030_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/spimemio/_0786_  (.A1(\soc/spimemio/_0168_ ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\soc/spimemio/_0157_ ),
    .C1(\soc/spimemio/_0321_ ),
    .C2(\soc/spimemio/_0214_ ),
    .Y(\soc/spimemio/_0031_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0788_  (.A1(\soc/spimemio/_0216_ ),
    .A2(\soc/spimemio/_0316_ ),
    .B1(\soc/spimemio/rd_addr[7] ),
    .Y(\soc/spimemio/_0330_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0789_  (.A(\soc/spimemio/rd_addr[7] ),
    .B(\soc/spimemio/_0216_ ),
    .Y(\soc/spimemio/_0331_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0790_  (.A1(net365),
    .A2(\soc/spimemio/_0309_ ),
    .B1(\soc/spimemio/_0317_ ),
    .B2(\soc/spimemio/_0331_ ),
    .Y(\soc/spimemio/_0332_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0791_  (.A1(\soc/spimemio/_0309_ ),
    .A2(\soc/spimemio/_0330_ ),
    .B1(\soc/spimemio/_0332_ ),
    .Y(\soc/spimemio/_0032_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0792_  (.A(\soc/spimemio/rd_inc ),
    .B(\soc/spimemio/_0181_ ),
    .Y(\soc/spimemio/_0333_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0793_  (.A(\soc/spimemio/_0316_ ),
    .B(\soc/spimemio/_0333_ ),
    .Y(\soc/spimemio/_0334_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0794_  (.A(\soc/spimemio/_0331_ ),
    .B(net106),
    .C(\soc/spimemio/_0333_ ),
    .Y(\soc/spimemio/_0335_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0795_  (.A1(net360),
    .A2(\soc/spimemio/_0306_ ),
    .B1(\soc/spimemio/_0334_ ),
    .B2(\soc/spimemio/rd_addr[8] ),
    .C1(\soc/spimemio/_0335_ ),
    .X(\soc/spimemio/_0033_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/spimemio/_0796_  (.A1(\soc/spimemio/_0178_ ),
    .A2(\soc/spimemio/_0181_ ),
    .A3(\soc/spimemio/_0317_ ),
    .B1(\soc/spimemio/_0309_ ),
    .B2(net355),
    .Y(\soc/spimemio/_0336_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0797_  (.A1(\soc/spimemio/_0178_ ),
    .A2(\soc/spimemio/_0334_ ),
    .B1(\soc/spimemio/_0336_ ),
    .Y(\soc/spimemio/_0034_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0798_  (.A(\soc/spimemio/_0212_ ),
    .B(\soc/spimemio/_0231_ ),
    .Y(\soc/spimemio/_0337_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0799_  (.A1(\soc/spimemio/rd_addr[10] ),
    .A2(\soc/spimemio/_0316_ ),
    .B1(\soc/spimemio/_0309_ ),
    .B2(net714),
    .Y(\soc/spimemio/_0338_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0800_  (.A1(\soc/spimemio/_0337_ ),
    .A2(\soc/spimemio/_0321_ ),
    .B1(net715),
    .Y(\soc/spimemio/_0035_ ));
 sky130_fd_sc_hd__nand4_1 \soc/spimemio/_0801_  (.A(\soc/spimemio/rd_addr[9] ),
    .B(\soc/spimemio/rd_addr[10] ),
    .C(\soc/spimemio/rd_addr[11] ),
    .D(\soc/spimemio/_0211_ ),
    .Y(\soc/spimemio/_0339_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/spimemio/_0802_  (.A1(\soc/spimemio/_0212_ ),
    .A2(net106),
    .B1(\soc/spimemio/_0309_ ),
    .C1(\soc/spimemio/_0179_ ),
    .Y(\soc/spimemio/_0340_ ));
 sky130_fd_sc_hd__o221a_1 \soc/spimemio/_0803_  (.A1(net744),
    .A2(\soc/spimemio/_0309_ ),
    .B1(\soc/spimemio/_0317_ ),
    .B2(\soc/spimemio/_0339_ ),
    .C1(\soc/spimemio/_0340_ ),
    .X(\soc/spimemio/_0036_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0804_  (.A(\iomem_addr[12] ),
    .B(\soc/spimemio/_0309_ ),
    .Y(\soc/spimemio/_0341_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0805_  (.A(\soc/spimemio/rd_addr[12] ),
    .B(\soc/spimemio/_0339_ ),
    .Y(\soc/spimemio/_0342_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_0806_  (.A1(\soc/spimemio/rd_addr[12] ),
    .A2(\soc/spimemio/_0316_ ),
    .B1(\soc/spimemio/_0317_ ),
    .B2(\soc/spimemio/_0342_ ),
    .Y(\soc/spimemio/_0343_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0807_  (.A(\soc/spimemio/_0341_ ),
    .B(\soc/spimemio/_0343_ ),
    .Y(\soc/spimemio/_0037_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0808_  (.A1(\soc/spimemio/rd_addr[12] ),
    .A2(\soc/spimemio/_0182_ ),
    .B1(\soc/spimemio/rd_addr[13] ),
    .Y(\soc/spimemio/_0344_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0809_  (.A1(\soc/spimemio/rd_addr[13] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[13] ),
    .Y(\soc/spimemio/_0345_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/spimemio/_0810_  (.A1(\soc/spimemio/_0206_ ),
    .A2(\soc/spimemio/_0317_ ),
    .A3(\soc/spimemio/_0344_ ),
    .B1(\soc/spimemio/_0345_ ),
    .Y(\soc/spimemio/_0038_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0811_  (.A(\soc/spimemio/rd_addr[14] ),
    .B(\soc/spimemio/_0206_ ),
    .Y(\soc/spimemio/_0346_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0812_  (.A(\soc/spimemio/_0183_ ),
    .B(\soc/spimemio/_0346_ ),
    .C(\soc/spimemio/_0317_ ),
    .Y(\soc/spimemio/_0347_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0813_  (.A1(\soc/spimemio/rd_addr[14] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(net947),
    .C1(\soc/spimemio/_0347_ ),
    .X(\soc/spimemio/_0039_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0814_  (.A1(\soc/spimemio/rd_addr[15] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[15] ),
    .Y(\soc/spimemio/_0348_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0815_  (.A1(\soc/spimemio/rd_addr[15] ),
    .A2(\soc/spimemio/_0183_ ),
    .B1(\soc/spimemio/_0317_ ),
    .Y(\soc/spimemio/_0349_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0816_  (.A1(\soc/spimemio/rd_addr[15] ),
    .A2(\soc/spimemio/_0183_ ),
    .B1(\soc/spimemio/_0349_ ),
    .Y(\soc/spimemio/_0350_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0817_  (.A(\soc/spimemio/_0348_ ),
    .B(\soc/spimemio/_0350_ ),
    .Y(\soc/spimemio/_0040_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0818_  (.A1(\soc/spimemio/rd_addr[15] ),
    .A2(\soc/spimemio/_0183_ ),
    .B1(\soc/spimemio/rd_addr[16] ),
    .Y(\soc/spimemio/_0351_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0819_  (.A(\soc/spimemio/_0202_ ),
    .B(\soc/spimemio/_0317_ ),
    .C(\soc/spimemio/_0351_ ),
    .Y(\soc/spimemio/_0352_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0820_  (.A1(\soc/spimemio/rd_addr[16] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[16] ),
    .C1(\soc/spimemio/_0352_ ),
    .X(\soc/spimemio/_0041_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0821_  (.A(\soc/spimemio/rd_addr[17] ),
    .B(\soc/spimemio/_0202_ ),
    .Y(\soc/spimemio/_0353_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0822_  (.A(\soc/spimemio/_0184_ ),
    .B(\soc/spimemio/_0317_ ),
    .C(\soc/spimemio/_0353_ ),
    .Y(\soc/spimemio/_0354_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0823_  (.A1(\soc/spimemio/rd_addr[17] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(net946),
    .C1(\soc/spimemio/_0354_ ),
    .X(\soc/spimemio/_0042_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0824_  (.A1(\soc/spimemio/rd_addr[18] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(net724),
    .Y(\soc/spimemio/_0355_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0825_  (.A1(\soc/spimemio/_0198_ ),
    .A2(\soc/spimemio/_0317_ ),
    .B1(\soc/spimemio/_0355_ ),
    .Y(\soc/spimemio/_0043_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0826_  (.A(\soc/spimemio/rd_addr[18] ),
    .B(\soc/spimemio/rd_addr[19] ),
    .C(\soc/spimemio/_0184_ ),
    .X(\soc/spimemio/_0356_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0827_  (.A1(\soc/spimemio/rd_addr[18] ),
    .A2(\soc/spimemio/_0184_ ),
    .B1(\soc/spimemio/rd_addr[19] ),
    .Y(\soc/spimemio/_0357_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0828_  (.A(\soc/spimemio/_0356_ ),
    .B(\soc/spimemio/_0317_ ),
    .C(\soc/spimemio/_0357_ ),
    .Y(\soc/spimemio/_0358_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0829_  (.A1(\soc/spimemio/rd_addr[19] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[19] ),
    .C1(\soc/spimemio/_0358_ ),
    .X(\soc/spimemio/_0044_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0830_  (.A(\soc/spimemio/rd_addr[20] ),
    .B(\soc/spimemio/_0356_ ),
    .Y(\soc/spimemio/_0359_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0831_  (.A(\soc/spimemio/_0186_ ),
    .B(\soc/spimemio/_0317_ ),
    .C(\soc/spimemio/_0359_ ),
    .Y(\soc/spimemio/_0360_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0832_  (.A1(\soc/spimemio/rd_addr[20] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[20] ),
    .C1(\soc/spimemio/_0360_ ),
    .X(\soc/spimemio/_0045_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0833_  (.A(\soc/spimemio/rd_addr[21] ),
    .B(\soc/spimemio/_0186_ ),
    .Y(\soc/spimemio/_0361_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0834_  (.A(\soc/spimemio/_0188_ ),
    .B(\soc/spimemio/_0317_ ),
    .C(\soc/spimemio/_0361_ ),
    .Y(\soc/spimemio/_0362_ ));
 sky130_fd_sc_hd__a221o_1 \soc/spimemio/_0835_  (.A1(\soc/spimemio/rd_addr[21] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[21] ),
    .C1(\soc/spimemio/_0362_ ),
    .X(\soc/spimemio/_0046_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/_0836_  (.A(\soc/spimemio/rd_addr[22] ),
    .B(\soc/spimemio/_0188_ ),
    .Y(\soc/spimemio/_0363_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0837_  (.A1(\soc/spimemio/rd_addr[22] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(\iomem_addr[22] ),
    .Y(\soc/spimemio/_0364_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0838_  (.A1(\soc/spimemio/_0363_ ),
    .A2(\soc/spimemio/_0317_ ),
    .B1(\soc/spimemio/_0364_ ),
    .Y(\soc/spimemio/_0047_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0839_  (.A(\soc/spimemio/_0192_ ),
    .B(\soc/spimemio/_0321_ ),
    .Y(\soc/spimemio/_0365_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0840_  (.A1(\soc/spimemio/rd_addr[23] ),
    .A2(net106),
    .B1(\soc/spimemio/_0306_ ),
    .B2(net694),
    .Y(\soc/spimemio/_0366_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0841_  (.A1(\soc/spimemio/_0190_ ),
    .A2(\soc/spimemio/_0365_ ),
    .B1(net695),
    .Y(\soc/spimemio/_0048_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0842_  (.A(net722),
    .B(\soc/spimemio/_0255_ ),
    .Y(\soc/spimemio/_0367_ ));
 sky130_fd_sc_hd__and4b_4 \soc/spimemio/_0843_  (.A_N(\soc/spimemio/dout_tag[3] ),
    .B(\soc/spimemio/_0367_ ),
    .C(\soc/spimemio/_0303_ ),
    .D(\soc/spimemio/dout_tag[1] ),
    .X(\soc/spimemio/_0368_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0845_  (.A0(\soc/spimemio/buffer[8] ),
    .A1(\soc/spimemio/dout_data[0] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0049_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0846_  (.A0(\soc/spimemio/buffer[9] ),
    .A1(\soc/spimemio/dout_data[1] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0050_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0847_  (.A0(\soc/spimemio/buffer[10] ),
    .A1(\soc/spimemio/dout_data[2] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0051_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0848_  (.A0(\soc/spimemio/buffer[11] ),
    .A1(\soc/spimemio/dout_data[3] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0052_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0849_  (.A0(\soc/spimemio/buffer[12] ),
    .A1(\soc/spimemio/dout_data[4] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0053_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0850_  (.A0(\soc/spimemio/buffer[13] ),
    .A1(\soc/spimemio/dout_data[5] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0054_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0851_  (.A0(\soc/spimemio/buffer[14] ),
    .A1(\soc/spimemio/dout_data[6] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0055_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0852_  (.A0(\soc/spimemio/buffer[15] ),
    .A1(\soc/spimemio/dout_data[7] ),
    .S(\soc/spimemio/_0368_ ),
    .X(\soc/spimemio/_0056_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0854_  (.A(\soc/spimemio/buffer[0] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0371_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0856_  (.A(\soc/spimem_rdata[0] ),
    .B(net107),
    .Y(\soc/spimemio/_0373_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0857_  (.A(\soc/spimemio/_0371_ ),
    .B(\soc/spimemio/_0373_ ),
    .Y(\soc/spimemio/_0057_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0858_  (.A(\soc/spimemio/buffer[1] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0374_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0859_  (.A(\soc/spimem_rdata[1] ),
    .B(\soc/spimemio/_0305_ ),
    .Y(\soc/spimemio/_0375_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0860_  (.A(\soc/spimemio/_0374_ ),
    .B(\soc/spimemio/_0375_ ),
    .Y(\soc/spimemio/_0058_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0861_  (.A(\soc/spimemio/buffer[2] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0376_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0862_  (.A(\soc/spimem_rdata[2] ),
    .B(net107),
    .Y(\soc/spimemio/_0377_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0863_  (.A(\soc/spimemio/_0376_ ),
    .B(\soc/spimemio/_0377_ ),
    .Y(\soc/spimemio/_0059_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0864_  (.A(\soc/spimemio/buffer[3] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0378_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0865_  (.A(\soc/spimem_rdata[3] ),
    .B(net107),
    .Y(\soc/spimemio/_0379_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0866_  (.A(\soc/spimemio/_0378_ ),
    .B(\soc/spimemio/_0379_ ),
    .Y(\soc/spimemio/_0060_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0867_  (.A(\soc/spimemio/buffer[4] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0380_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0868_  (.A(\soc/spimem_rdata[4] ),
    .B(net107),
    .Y(\soc/spimemio/_0381_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0869_  (.A(\soc/spimemio/_0380_ ),
    .B(\soc/spimemio/_0381_ ),
    .Y(\soc/spimemio/_0061_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0870_  (.A(\soc/spimemio/buffer[5] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0382_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0871_  (.A(\soc/spimem_rdata[5] ),
    .B(net107),
    .Y(\soc/spimemio/_0383_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0872_  (.A(\soc/spimemio/_0382_ ),
    .B(\soc/spimemio/_0383_ ),
    .Y(\soc/spimemio/_0062_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0873_  (.A(\soc/spimemio/buffer[6] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0384_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0874_  (.A(\soc/spimem_rdata[6] ),
    .B(\soc/spimemio/_0305_ ),
    .Y(\soc/spimemio/_0385_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0875_  (.A(\soc/spimemio/_0384_ ),
    .B(\soc/spimemio/_0385_ ),
    .Y(\soc/spimemio/_0063_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0876_  (.A(\soc/spimemio/buffer[7] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0386_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0877_  (.A(\soc/spimem_rdata[7] ),
    .B(net107),
    .Y(\soc/spimemio/_0387_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0878_  (.A(\soc/spimemio/_0386_ ),
    .B(\soc/spimemio/_0387_ ),
    .Y(\soc/spimemio/_0064_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0879_  (.A(\soc/spimemio/buffer[8] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0388_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0880_  (.A(\soc/spimem_rdata[8] ),
    .B(net107),
    .Y(\soc/spimemio/_0389_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0881_  (.A(\soc/spimemio/_0388_ ),
    .B(\soc/spimemio/_0389_ ),
    .Y(\soc/spimemio/_0065_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0882_  (.A(\soc/spimemio/buffer[9] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0390_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0883_  (.A(\soc/spimem_rdata[9] ),
    .B(net107),
    .Y(\soc/spimemio/_0391_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0884_  (.A(\soc/spimemio/_0390_ ),
    .B(\soc/spimemio/_0391_ ),
    .Y(\soc/spimemio/_0066_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0886_  (.A(\soc/spimemio/buffer[10] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0393_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0888_  (.A(\soc/spimem_rdata[10] ),
    .B(net107),
    .Y(\soc/spimemio/_0395_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0889_  (.A(\soc/spimemio/_0393_ ),
    .B(\soc/spimemio/_0395_ ),
    .Y(\soc/spimemio/_0067_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0890_  (.A(net710),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0396_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0891_  (.A(\soc/spimem_rdata[11] ),
    .B(net107),
    .Y(\soc/spimemio/_0397_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0892_  (.A(net711),
    .B(\soc/spimemio/_0397_ ),
    .Y(\soc/spimemio/_0068_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0893_  (.A(\soc/spimemio/buffer[12] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0398_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0894_  (.A(\soc/spimem_rdata[12] ),
    .B(net107),
    .Y(\soc/spimemio/_0399_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0895_  (.A(\soc/spimemio/_0398_ ),
    .B(\soc/spimemio/_0399_ ),
    .Y(\soc/spimemio/_0069_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0896_  (.A(\soc/spimemio/buffer[13] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0400_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0897_  (.A(\soc/spimem_rdata[13] ),
    .B(net107),
    .Y(\soc/spimemio/_0401_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0898_  (.A(\soc/spimemio/_0400_ ),
    .B(\soc/spimemio/_0401_ ),
    .Y(\soc/spimemio/_0070_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0899_  (.A(\soc/spimemio/buffer[14] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0402_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0900_  (.A(\soc/spimem_rdata[14] ),
    .B(net107),
    .Y(\soc/spimemio/_0403_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0901_  (.A(\soc/spimemio/_0402_ ),
    .B(\soc/spimemio/_0403_ ),
    .Y(\soc/spimemio/_0071_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0902_  (.A(\soc/spimemio/buffer[15] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0404_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0903_  (.A(\soc/spimem_rdata[15] ),
    .B(net107),
    .Y(\soc/spimemio/_0405_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0904_  (.A(\soc/spimemio/_0404_ ),
    .B(\soc/spimemio/_0405_ ),
    .Y(\soc/spimemio/_0072_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0905_  (.A(\soc/spimemio/buffer[16] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0406_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0906_  (.A(\soc/spimem_rdata[16] ),
    .B(net107),
    .Y(\soc/spimemio/_0407_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0907_  (.A(\soc/spimemio/_0406_ ),
    .B(\soc/spimemio/_0407_ ),
    .Y(\soc/spimemio/_0073_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0908_  (.A(\soc/spimemio/buffer[17] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0408_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0909_  (.A(\soc/spimem_rdata[17] ),
    .B(net107),
    .Y(\soc/spimemio/_0409_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0910_  (.A(\soc/spimemio/_0408_ ),
    .B(\soc/spimemio/_0409_ ),
    .Y(\soc/spimemio/_0074_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0911_  (.A(\soc/spimemio/buffer[18] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0410_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0912_  (.A(\soc/spimem_rdata[18] ),
    .B(net106),
    .Y(\soc/spimemio/_0411_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0913_  (.A(\soc/spimemio/_0410_ ),
    .B(\soc/spimemio/_0411_ ),
    .Y(\soc/spimemio/_0075_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0914_  (.A(\soc/spimemio/buffer[19] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0412_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0915_  (.A(\soc/spimem_rdata[19] ),
    .B(net107),
    .Y(\soc/spimemio/_0413_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0916_  (.A(\soc/spimemio/_0412_ ),
    .B(\soc/spimemio/_0413_ ),
    .Y(\soc/spimemio/_0076_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0918_  (.A(net841),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0415_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0920_  (.A(\soc/spimem_rdata[20] ),
    .B(net107),
    .Y(\soc/spimemio/_0417_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0921_  (.A(\soc/spimemio/_0415_ ),
    .B(\soc/spimemio/_0417_ ),
    .Y(\soc/spimemio/_0077_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0922_  (.A(\soc/spimemio/buffer[21] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0418_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0923_  (.A(\soc/spimem_rdata[21] ),
    .B(net107),
    .Y(\soc/spimemio/_0419_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0924_  (.A(\soc/spimemio/_0418_ ),
    .B(\soc/spimemio/_0419_ ),
    .Y(\soc/spimemio/_0078_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0925_  (.A(\soc/spimemio/buffer[22] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0420_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0926_  (.A(\soc/spimem_rdata[22] ),
    .B(net106),
    .Y(\soc/spimemio/_0421_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0927_  (.A(\soc/spimemio/_0420_ ),
    .B(\soc/spimemio/_0421_ ),
    .Y(\soc/spimemio/_0079_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0928_  (.A(\soc/spimemio/buffer[23] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0422_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0929_  (.A(\soc/spimem_rdata[23] ),
    .B(net107),
    .Y(\soc/spimemio/_0423_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0930_  (.A(\soc/spimemio/_0422_ ),
    .B(\soc/spimemio/_0423_ ),
    .Y(\soc/spimemio/_0080_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0931_  (.A(\soc/spimemio/dout_data[0] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0424_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0932_  (.A(\soc/spimem_rdata[24] ),
    .B(net107),
    .Y(\soc/spimemio/_0425_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0933_  (.A(\soc/spimemio/_0424_ ),
    .B(\soc/spimemio/_0425_ ),
    .Y(\soc/spimemio/_0081_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0934_  (.A(\soc/spimemio/dout_data[1] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0426_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0935_  (.A(\soc/spimem_rdata[25] ),
    .B(net107),
    .Y(\soc/spimemio/_0427_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0936_  (.A(\soc/spimemio/_0426_ ),
    .B(\soc/spimemio/_0427_ ),
    .Y(\soc/spimemio/_0082_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0937_  (.A(\soc/spimemio/dout_data[2] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0428_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0938_  (.A(\soc/spimem_rdata[26] ),
    .B(net106),
    .Y(\soc/spimemio/_0429_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0939_  (.A(\soc/spimemio/_0428_ ),
    .B(\soc/spimemio/_0429_ ),
    .Y(\soc/spimemio/_0083_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0940_  (.A(\soc/spimemio/dout_data[3] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0430_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0941_  (.A(\soc/spimem_rdata[27] ),
    .B(net107),
    .Y(\soc/spimemio/_0431_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0942_  (.A(\soc/spimemio/_0430_ ),
    .B(\soc/spimemio/_0431_ ),
    .Y(\soc/spimemio/_0084_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0943_  (.A(\soc/spimemio/dout_data[4] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0432_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0944_  (.A(\soc/spimem_rdata[28] ),
    .B(net107),
    .Y(\soc/spimemio/_0433_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0945_  (.A(\soc/spimemio/_0432_ ),
    .B(\soc/spimemio/_0433_ ),
    .Y(\soc/spimemio/_0085_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0946_  (.A(\soc/spimemio/dout_data[5] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0434_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0947_  (.A(\soc/spimem_rdata[29] ),
    .B(net107),
    .Y(\soc/spimemio/_0435_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0948_  (.A(\soc/spimemio/_0434_ ),
    .B(\soc/spimemio/_0435_ ),
    .Y(\soc/spimemio/_0086_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0949_  (.A(\soc/spimemio/dout_data[6] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0436_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0950_  (.A(\soc/spimem_rdata[30] ),
    .B(net107),
    .Y(\soc/spimemio/_0437_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0951_  (.A(\soc/spimemio/_0436_ ),
    .B(\soc/spimemio/_0437_ ),
    .Y(\soc/spimemio/_0087_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0952_  (.A(\soc/spimemio/dout_data[7] ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0438_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0953_  (.A(\soc/spimem_rdata[31] ),
    .B(net107),
    .Y(\soc/spimemio/_0439_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0954_  (.A(\soc/spimemio/_0438_ ),
    .B(\soc/spimemio/_0439_ ),
    .Y(\soc/spimemio/_0088_ ));
 sky130_fd_sc_hd__or3_1 \soc/spimemio/_0955_  (.A(\soc/spimemio/state[6] ),
    .B(\soc/spimemio/state[5] ),
    .C(\soc/spimemio/state[12] ),
    .X(\soc/spimemio/_0440_ ));
 sky130_fd_sc_hd__or3_1 \soc/spimemio/_0956_  (.A(\soc/spimemio/state[4] ),
    .B(\soc/spimemio/state[2] ),
    .C(\soc/spimemio/state[1] ),
    .X(\soc/spimemio/_0441_ ));
 sky130_fd_sc_hd__or3_2 \soc/spimemio/_0957_  (.A(\soc/spimemio/state[9] ),
    .B(\soc/spimemio/_0440_ ),
    .C(\soc/spimemio/_0441_ ),
    .X(\soc/spimemio/_0442_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0958_  (.A(\soc/spimemio/state[0] ),
    .B(\soc/spimemio/_0442_ ),
    .Y(\soc/spimemio/_0443_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0959_  (.A(\soc/spimemio/_0245_ ),
    .B(\soc/spimemio/_0280_ ),
    .Y(\soc/spimemio/_0444_ ));
 sky130_fd_sc_hd__nor2_4 \soc/spimemio/_0960_  (.A(\soc/spimemio/_0443_ ),
    .B(\soc/spimemio/_0444_ ),
    .Y(\soc/spimemio/_0445_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0961_  (.A1(\soc/spimemio/_0273_ ),
    .A2(\soc/spimemio_cfgreg_do[16] ),
    .B1(\soc/spimemio/state[1] ),
    .Y(\soc/spimemio/_0446_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/spimemio/_0962_  (.A1(net736),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[6] ),
    .B2(net362),
    .C1(net456),
    .C2(\soc/spimemio/_0277_ ),
    .Y(\soc/spimemio/_0447_ ));
 sky130_fd_sc_hd__and4_1 \soc/spimemio/_0963_  (.A(\soc/spimemio/_0263_ ),
    .B(\soc/spimemio/_0269_ ),
    .C(\soc/spimemio/_0446_ ),
    .D(\soc/spimemio/_0447_ ),
    .X(\soc/spimemio/_0448_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0965_  (.A(\soc/spimemio/din_data[0] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0450_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_0966_  (.A1(\soc/spimemio/_0442_ ),
    .A2(\soc/spimemio/_0445_ ),
    .A3(net737),
    .B1(\soc/spimemio/_0450_ ),
    .Y(\soc/spimemio/_0091_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/spimemio/_0967_  (.A1(\soc/spimemio/config_cont ),
    .A2(\soc/spimemio/_0274_ ),
    .B1(\soc/spimemio/_0442_ ),
    .Y(\soc/spimemio/_0451_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0968_  (.A(\soc/spimemio/xfer/_047_ ),
    .B(\soc/spimemio/state[1] ),
    .C(\soc/spimemio_cfgreg_do[17] ),
    .Y(\soc/spimemio/_0452_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0969_  (.A1(net356),
    .A2(\soc/spimemio/state[6] ),
    .B1(\soc/spimemio/state[4] ),
    .Y(\soc/spimemio/_0453_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0970_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/config_qspi ),
    .Y(\soc/spimemio/_0454_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/spimemio/_0971_  (.A1(net779),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[2] ),
    .B2(\soc/spimemio/_0454_ ),
    .C1(\soc/spimemio/_0277_ ),
    .C2(net457),
    .Y(\soc/spimemio/_0455_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0972_  (.A(\soc/spimemio/_0452_ ),
    .B(\soc/spimemio/_0453_ ),
    .C(\soc/spimemio/_0455_ ),
    .Y(\soc/spimemio/_0456_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0973_  (.A(\soc/spimemio/_0451_ ),
    .B(\soc/spimemio/_0456_ ),
    .Y(\soc/spimemio/_0457_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0974_  (.A(\soc/spimemio/din_data[1] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0458_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0975_  (.A1(\soc/spimemio/_0445_ ),
    .A2(\soc/spimemio/_0457_ ),
    .B1(\soc/spimemio/_0458_ ),
    .Y(\soc/spimemio/_0092_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/spimemio/_0976_  (.A1(net724),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[1] ),
    .B2(\soc/spimemio_cfgreg_do[18] ),
    .C1(\soc/spimemio/_0277_ ),
    .C2(net394),
    .Y(\soc/spimemio/_0459_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0977_  (.A(net714),
    .B(\soc/spimemio/state[6] ),
    .Y(\soc/spimemio/_0460_ ));
 sky130_fd_sc_hd__o211a_1 \soc/spimemio/_0978_  (.A1(\soc/spimemio/_0269_ ),
    .A2(\soc/spimemio/_0454_ ),
    .B1(\soc/spimemio/_0460_ ),
    .C1(\soc/spimemio/_0274_ ),
    .X(\soc/spimemio/_0461_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0979_  (.A(\soc/spimemio/_0442_ ),
    .B(\soc/spimemio/_0459_ ),
    .C(\soc/spimemio/_0461_ ),
    .Y(\soc/spimemio/_0462_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_0980_  (.A0(\soc/spimemio/din_data[2] ),
    .A1(\soc/spimemio/_0462_ ),
    .S(\soc/spimemio/_0445_ ),
    .X(\soc/spimemio/_0093_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0981_  (.A1(\iomem_addr[19] ),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[6] ),
    .B2(net744),
    .Y(\soc/spimemio/_0463_ ));
 sky130_fd_sc_hd__o21ai_1 \soc/spimemio/_0982_  (.A1(\soc/spimemio/config_ddr ),
    .A2(\soc/spimemio/config_qspi ),
    .B1(\soc/spimemio/state[2] ),
    .Y(\soc/spimemio/_0464_ ));
 sky130_fd_sc_hd__a32oi_1 \soc/spimemio/_0983_  (.A1(\soc/spimemio/xfer/_047_ ),
    .A2(\soc/spimemio/state[1] ),
    .A3(net756),
    .B1(\soc/spimemio/_0277_ ),
    .B2(net387),
    .Y(\soc/spimemio/_0465_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_0984_  (.A(\soc/spimemio/_0463_ ),
    .B(\soc/spimemio/_0464_ ),
    .C(\soc/spimemio/_0465_ ),
    .Y(\soc/spimemio/_0466_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_0985_  (.A(\soc/spimemio/state[4] ),
    .B(\soc/spimemio/_0451_ ),
    .C(\soc/spimemio/_0466_ ),
    .Y(\soc/spimemio/_0467_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0986_  (.A(\soc/spimemio/din_data[3] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0468_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0987_  (.A1(\soc/spimemio/_0445_ ),
    .A2(\soc/spimemio/_0467_ ),
    .B1(\soc/spimemio/_0468_ ),
    .Y(\soc/spimemio/_0094_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0988_  (.A(\soc/spimemio/state[2] ),
    .B(\soc/spimemio/config_ddr ),
    .Y(\soc/spimemio/_0469_ ));
 sky130_fd_sc_hd__a222oi_1 \soc/spimemio/_0989_  (.A1(\iomem_addr[20] ),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[6] ),
    .B2(net771),
    .C1(net381),
    .C2(\soc/spimemio/_0277_ ),
    .Y(\soc/spimemio/_0470_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_0990_  (.A1(\soc/spimemio/config_qspi ),
    .A2(\soc/spimemio/_0469_ ),
    .B1(\soc/spimemio/_0470_ ),
    .Y(\soc/spimemio/_0471_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0991_  (.A(\soc/spimemio/_0451_ ),
    .B(\soc/spimemio/_0471_ ),
    .Y(\soc/spimemio/_0472_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0992_  (.A(\soc/spimemio/din_data[4] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0473_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0993_  (.A1(\soc/spimemio/_0445_ ),
    .A2(\soc/spimemio/_0472_ ),
    .B1(\soc/spimemio/_0473_ ),
    .Y(\soc/spimemio/_0095_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_0994_  (.A(\soc/spimemio/_0263_ ),
    .B(\soc/spimemio/_0274_ ),
    .C(\soc/spimemio/_0442_ ),
    .X(\soc/spimemio/_0474_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_0995_  (.A1(\iomem_addr[21] ),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[6] ),
    .B2(\iomem_addr[13] ),
    .Y(\soc/spimemio/_0475_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_0996_  (.A(\soc/spimemio/_0464_ ),
    .B(\soc/spimemio/_0475_ ),
    .Y(\soc/spimemio/_0476_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_0997_  (.A1(net374),
    .A2(\soc/spimemio/_0277_ ),
    .B1(\soc/spimemio/_0476_ ),
    .Y(\soc/spimemio/_0477_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_0998_  (.A(\soc/spimemio/din_data[5] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0478_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_0999_  (.A1(\soc/spimemio/_0445_ ),
    .A2(\soc/spimemio/_0474_ ),
    .A3(\soc/spimemio/_0477_ ),
    .B1(\soc/spimemio/_0478_ ),
    .Y(\soc/spimemio/_0096_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_1000_  (.A1(\soc/spimemio/state[2] ),
    .A2(\soc/spimemio/config_qspi ),
    .B1(\soc/spimemio/_0277_ ),
    .B2(net505),
    .Y(\soc/spimemio/_0479_ ));
 sky130_fd_sc_hd__a221oi_1 \soc/spimemio/_1001_  (.A1(\iomem_addr[22] ),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[6] ),
    .B2(net708),
    .C1(\soc/spimemio/_0451_ ),
    .Y(\soc/spimemio/_0480_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1002_  (.A(\soc/spimemio/din_data[6] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0481_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_1003_  (.A1(\soc/spimemio/_0445_ ),
    .A2(\soc/spimemio/_0479_ ),
    .A3(net709),
    .B1(\soc/spimemio/_0481_ ),
    .Y(\soc/spimemio/_0097_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/_1004_  (.A1(net694),
    .A2(\soc/spimemio/state[9] ),
    .B1(\soc/spimemio/state[6] ),
    .B2(net713),
    .Y(\soc/spimemio/_0482_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1005_  (.A(\soc/spimemio/_0464_ ),
    .B(\soc/spimemio/_0482_ ),
    .Y(\soc/spimemio/_0483_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_1006_  (.A1(net365),
    .A2(\soc/spimemio/_0277_ ),
    .B1(\soc/spimemio/_0483_ ),
    .Y(\soc/spimemio/_0484_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1007_  (.A(\soc/spimemio/din_data[7] ),
    .B(\soc/spimemio/_0445_ ),
    .Y(\soc/spimemio/_0485_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_1008_  (.A1(\soc/spimemio/_0445_ ),
    .A2(\soc/spimemio/_0474_ ),
    .A3(\soc/spimemio/_0484_ ),
    .B1(\soc/spimemio/_0485_ ),
    .Y(\soc/spimemio/_0098_ ));
 sky130_fd_sc_hd__nand4_4 \soc/spimemio/_1009_  (.A(\soc/spimemio/dout_tag[0] ),
    .B(\soc/spimemio/dout_valid ),
    .C(\soc/spimemio/_0367_ ),
    .D(\soc/spimemio/_0304_ ),
    .Y(\soc/spimemio/_0486_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1010_  (.A0(\soc/spimemio/dout_data[0] ),
    .A1(\soc/spimemio/buffer[0] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0102_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1011_  (.A0(\soc/spimemio/dout_data[1] ),
    .A1(\soc/spimemio/buffer[1] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0103_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1012_  (.A0(\soc/spimemio/dout_data[2] ),
    .A1(\soc/spimemio/buffer[2] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0104_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1013_  (.A0(\soc/spimemio/dout_data[3] ),
    .A1(\soc/spimemio/buffer[3] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0105_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1014_  (.A0(\soc/spimemio/dout_data[4] ),
    .A1(\soc/spimemio/buffer[4] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0106_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1015_  (.A0(\soc/spimemio/dout_data[5] ),
    .A1(\soc/spimemio/buffer[5] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0107_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1016_  (.A0(\soc/spimemio/dout_data[6] ),
    .A1(\soc/spimemio/buffer[6] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0108_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/_1017_  (.A0(\soc/spimemio/dout_data[7] ),
    .A1(\soc/spimemio/buffer[7] ),
    .S(\soc/spimemio/_0486_ ),
    .X(\soc/spimemio/_0109_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1018_  (.A1(\soc/spimemio/rd_wait ),
    .A2(\soc/spimemio/_0316_ ),
    .B1(\soc/spimemio/_0309_ ),
    .Y(\soc/spimemio/_0487_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_1019_  (.A1(net727),
    .A2(\soc/spimemio/_0245_ ),
    .B1(\soc/spimemio/_0487_ ),
    .Y(\soc/spimemio/_0111_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1020_  (.A(\soc/spimemio/rd_inc ),
    .B(\soc/spimemio/_0316_ ),
    .Y(\soc/spimemio/_0488_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_1021_  (.A1(\soc/spimemio/_0269_ ),
    .A2(net733),
    .B1(\soc/spimemio/_0255_ ),
    .Y(\soc/spimemio/_0489_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1022_  (.A(\soc/spimemio/_0488_ ),
    .B(\soc/spimemio/_0489_ ),
    .Y(\soc/spimemio/_0112_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1023_  (.A1(\soc/spimemio/state[7] ),
    .A2(\soc/spimemio/state[10] ),
    .B1(\soc/spimemio/dout_valid ),
    .Y(\soc/spimemio/_0490_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/_1024_  (.A(net733),
    .B(\soc/spimemio/_0245_ ),
    .C(\soc/spimemio/_0490_ ),
    .X(\soc/spimemio/_0089_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_1025_  (.A1(\soc/spimemio/xfer/_047_ ),
    .A2(\soc/spimemio/state[1] ),
    .B1(\soc/spimemio/din_rd ),
    .Y(\soc/spimemio/_0491_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1026_  (.A(\soc/spimemio/_0246_ ),
    .B(\soc/spimemio/_0491_ ),
    .Y(\soc/spimemio/_0100_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_1027_  (.A1(\soc/spimemio/_0241_ ),
    .A2(\soc/spimemio/_0315_ ),
    .B1(\soc/spimemio/_0246_ ),
    .Y(\soc/spimemio/_0110_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1028_  (.A(\soc/spimemio/state[9] ),
    .B(\soc/spimemio/state[3] ),
    .Y(\soc/spimemio/_0492_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1029_  (.A(\soc/spimemio/_0259_ ),
    .B(\soc/spimemio/_0264_ ),
    .Y(\soc/spimemio/_0493_ ));
 sky130_fd_sc_hd__nor4_1 \soc/spimemio/_1030_  (.A(\soc/spimemio/state[0] ),
    .B(\soc/spimemio/_0440_ ),
    .C(\soc/spimemio/_0441_ ),
    .D(\soc/spimemio/_0493_ ),
    .Y(\soc/spimemio/_0494_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1031_  (.A(\soc/spimemio/_0265_ ),
    .B(\soc/spimemio/_0280_ ),
    .Y(\soc/spimemio/_0495_ ));
 sky130_fd_sc_hd__a21oi_2 \soc/spimemio/_1032_  (.A1(\soc/spimemio/_0492_ ),
    .A2(\soc/spimemio/_0494_ ),
    .B1(\soc/spimemio/_0495_ ),
    .Y(\soc/spimemio/_0496_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1033_  (.A1(\soc/spimemio/din_tag[0] ),
    .A2(\soc/spimemio/_0496_ ),
    .B1(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0497_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_1034_  (.A1(\soc/spimemio/_0259_ ),
    .A2(\soc/spimemio/_0264_ ),
    .A3(\soc/spimemio/_0496_ ),
    .B1(\soc/spimemio/_0497_ ),
    .Y(\soc/spimemio/_0022_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1035_  (.A1(\soc/spimemio/din_tag[1] ),
    .A2(\soc/spimemio/_0496_ ),
    .B1(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0498_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/_1036_  (.A1(\soc/spimemio/_0261_ ),
    .A2(\soc/spimemio/_0264_ ),
    .A3(\soc/spimemio/_0496_ ),
    .B1(\soc/spimemio/_0498_ ),
    .Y(\soc/spimemio/_0023_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1037_  (.A(\soc/spimemio/state[3] ),
    .B(\soc/spimemio/_0266_ ),
    .Y(\soc/spimemio/_0499_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1038_  (.A(\soc/spimemio/din_tag[2] ),
    .B(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0500_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/_1039_  (.A1(\soc/spimemio/_0499_ ),
    .A2(\soc/spimemio/_0444_ ),
    .B1(\soc/spimemio/_0496_ ),
    .B2(\soc/spimemio/_0500_ ),
    .Y(\soc/spimemio/_0024_ ));
 sky130_fd_sc_hd__o211ai_2 \soc/spimemio/_1040_  (.A1(\soc/spimemio/_0242_ ),
    .A2(\soc/spimemio/_0492_ ),
    .B1(\soc/spimemio/_0494_ ),
    .C1(\soc/spimemio/_0499_ ),
    .Y(\soc/spimemio/_0501_ ));
 sky130_fd_sc_hd__and2_0 \soc/spimemio/_1041_  (.A(\soc/spimemio/_0257_ ),
    .B(\soc/spimemio/_0501_ ),
    .X(\soc/spimemio/_0090_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1042_  (.A(\soc/spimemio/config_cont ),
    .B(\soc/spimemio/_0244_ ),
    .Y(\soc/spimemio/_0502_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1043_  (.A(\soc/spimemio/din_qspi ),
    .B(\soc/spimemio/_0251_ ),
    .Y(\soc/spimemio/_0503_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1044_  (.A1(\soc/spimemio/config_qspi ),
    .A2(\soc/spimemio/_0252_ ),
    .B1(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0504_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_1045_  (.A(\soc/spimemio/_0502_ ),
    .B(\soc/spimemio/_0503_ ),
    .C(\soc/spimemio/_0504_ ),
    .Y(\soc/spimemio/_0099_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1046_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/spimemio/_0252_ ),
    .Y(\soc/spimemio/_0505_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1047_  (.A1(\soc/spimemio/din_ddr ),
    .A2(\soc/spimemio/_0251_ ),
    .B1(\soc/spimemio/_0245_ ),
    .Y(\soc/spimemio/_0506_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_1048_  (.A(\soc/spimemio/_0502_ ),
    .B(\soc/spimemio/_0505_ ),
    .C(\soc/spimemio/_0506_ ),
    .Y(\soc/spimemio/_0101_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/_1051_  (.A_N(\soc/_007_ ),
    .B(\soc/spimemio/config_en ),
    .Y(\soc/spimemio/_0509_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1052_  (.A(\soc/_007_ ),
    .B(net165),
    .Y(\soc/spimemio/_0510_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/_1053_  (.A(_074_),
    .B(\soc/spimemio/_0509_ ),
    .C(\soc/spimemio/_0510_ ),
    .Y(\soc/spimemio/_0113_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1054_  (.A(\soc/spimemio/config_ddr ),
    .B(\soc/_006_ ),
    .Y(\soc/spimemio/_0511_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_1055_  (.A(\soc/_006_ ),
    .Y(\soc/spimemio/_0512_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1056_  (.A1(\soc/spimemio/_0512_ ),
    .A2(net192),
    .B1(_074_),
    .Y(\soc/spimemio/_0513_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1057_  (.A(\soc/spimemio/_0511_ ),
    .B(\soc/spimemio/_0513_ ),
    .Y(\soc/spimemio/_0114_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1058_  (.A(\soc/spimemio/config_qspi ),
    .B(\soc/_006_ ),
    .Y(\soc/spimemio/_0514_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1059_  (.A1(\soc/spimemio/_0512_ ),
    .A2(net195),
    .B1(_074_),
    .Y(\soc/spimemio/_0515_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1060_  (.A(\soc/spimemio/_0514_ ),
    .B(\soc/spimemio/_0515_ ),
    .Y(\soc/spimemio/_0115_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1061_  (.A1(\soc/spimemio/_0512_ ),
    .A2(net199),
    .B1(_074_),
    .Y(\soc/spimemio/_0516_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/_1062_  (.A1(\soc/spimemio/_0279_ ),
    .A2(\soc/spimemio/_0512_ ),
    .B1(\soc/spimemio/_0516_ ),
    .Y(\soc/spimemio/_0116_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1063_  (.A(\soc/_006_ ),
    .B(\soc/spimemio_cfgreg_do[16] ),
    .Y(\soc/spimemio/_0517_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1064_  (.A1(\soc/spimemio/_0512_ ),
    .A2(net212),
    .B1(_074_),
    .Y(\soc/spimemio/_0518_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1065_  (.A(\soc/spimemio/_0517_ ),
    .B(\soc/spimemio/_0518_ ),
    .Y(\soc/spimemio/_0117_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1066_  (.A(\soc/_006_ ),
    .B(\soc/spimemio_cfgreg_do[17] ),
    .Y(\soc/spimemio/_0519_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1067_  (.A1(\soc/spimemio/_0512_ ),
    .A2(net209),
    .B1(_074_),
    .Y(\soc/spimemio/_0520_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1068_  (.A(\soc/spimemio/_0519_ ),
    .B(\soc/spimemio/_0520_ ),
    .Y(\soc/spimemio/_0118_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1069_  (.A(\soc/_006_ ),
    .B(\soc/spimemio_cfgreg_do[18] ),
    .Y(\soc/spimemio/_0521_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1070_  (.A1(\soc/spimemio/_0512_ ),
    .A2(net206),
    .B1(_074_),
    .Y(\soc/spimemio/_0522_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1071_  (.A(\soc/spimemio/_0521_ ),
    .B(\soc/spimemio/_0522_ ),
    .Y(\soc/spimemio/_0119_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/spimemio/_1072_  (.A0(\soc/spimemio_cfgreg_do[19] ),
    .A1(net202),
    .S(\soc/_006_ ),
    .Y(\soc/spimemio/_0523_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/_1073_  (.A(_074_),
    .B(\soc/spimemio/_0523_ ),
    .Y(\soc/spimemio/_0120_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1074_  (.A(\soc/_005_ ),
    .B(\soc/spimemio/config_oe[0] ),
    .Y(\soc/spimemio/_0524_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_1075_  (.A(\soc/_005_ ),
    .Y(\soc/spimemio/_0525_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1076_  (.A1(\soc/spimemio/_0525_ ),
    .A2(net244),
    .B1(_074_),
    .Y(\soc/spimemio/_0526_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1077_  (.A(\soc/spimemio/_0524_ ),
    .B(\soc/spimemio/_0526_ ),
    .Y(\soc/spimemio/_0121_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1078_  (.A(\soc/_005_ ),
    .B(\soc/spimemio/config_oe[1] ),
    .Y(\soc/spimemio/_0527_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1079_  (.A1(\soc/spimemio/_0525_ ),
    .A2(net237),
    .B1(_074_),
    .Y(\soc/spimemio/_0528_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1080_  (.A(\soc/spimemio/_0527_ ),
    .B(\soc/spimemio/_0528_ ),
    .Y(\soc/spimemio/_0122_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1081_  (.A(\soc/_005_ ),
    .B(\soc/spimemio/config_oe[2] ),
    .Y(\soc/spimemio/_0529_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1082_  (.A1(\soc/spimemio/_0525_ ),
    .A2(net235),
    .B1(_074_),
    .Y(\soc/spimemio/_0530_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1083_  (.A(\soc/spimemio/_0529_ ),
    .B(\soc/spimemio/_0530_ ),
    .Y(\soc/spimemio/_0123_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1084_  (.A(\soc/_005_ ),
    .B(\soc/spimemio/config_oe[3] ),
    .Y(\soc/spimemio/_0531_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1085_  (.A1(\soc/spimemio/_0525_ ),
    .A2(net231),
    .B1(_074_),
    .Y(\soc/spimemio/_0532_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1086_  (.A(\soc/spimemio/_0531_ ),
    .B(\soc/spimemio/_0532_ ),
    .Y(\soc/spimemio/_0124_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1087_  (.A(\soc/_004_ ),
    .B(\soc/spimemio/config_csb ),
    .Y(\soc/spimemio/_0533_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_1088_  (.A(\soc/_004_ ),
    .Y(\soc/spimemio/_0534_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1089_  (.A1(\soc/spimemio/_0534_ ),
    .A2(net263),
    .B1(_074_),
    .Y(\soc/spimemio/_0535_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1090_  (.A(\soc/spimemio/_0533_ ),
    .B(\soc/spimemio/_0535_ ),
    .Y(\soc/spimemio/_0125_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1091_  (.A(\soc/_004_ ),
    .B(\soc/spimemio/config_clk ),
    .Y(\soc/spimemio/_0536_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1092_  (.A1(\soc/spimemio/_0534_ ),
    .A2(net265),
    .B1(_074_),
    .Y(\soc/spimemio/_0537_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1093_  (.A(\soc/spimemio/_0536_ ),
    .B(\soc/spimemio/_0537_ ),
    .Y(\soc/spimemio/_0126_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1094_  (.A(\soc/_004_ ),
    .B(\soc/spimemio/config_do[0] ),
    .Y(\soc/spimemio/_0538_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1095_  (.A1(\soc/spimemio/_0534_ ),
    .A2(net286),
    .B1(_074_),
    .Y(\soc/spimemio/_0539_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1096_  (.A(\soc/spimemio/_0538_ ),
    .B(\soc/spimemio/_0539_ ),
    .Y(\soc/spimemio/_0127_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1097_  (.A(\soc/_004_ ),
    .B(\soc/spimemio/config_do[1] ),
    .Y(\soc/spimemio/_0540_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1098_  (.A1(\soc/spimemio/_0534_ ),
    .A2(net279),
    .B1(_074_),
    .Y(\soc/spimemio/_0541_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1099_  (.A(\soc/spimemio/_0540_ ),
    .B(\soc/spimemio/_0541_ ),
    .Y(\soc/spimemio/_0128_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1100_  (.A(\soc/_004_ ),
    .B(\soc/spimemio/config_do[2] ),
    .Y(\soc/spimemio/_0542_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1101_  (.A1(\soc/spimemio/_0534_ ),
    .A2(net271),
    .B1(_074_),
    .Y(\soc/spimemio/_0543_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1102_  (.A(\soc/spimemio/_0542_ ),
    .B(\soc/spimemio/_0543_ ),
    .Y(\soc/spimemio/_0129_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1103_  (.A(\soc/_004_ ),
    .B(\soc/spimemio/config_do[3] ),
    .Y(\soc/spimemio/_0544_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/_1104_  (.A1(\soc/spimemio/_0534_ ),
    .A2(net267),
    .B1(_074_),
    .Y(\soc/spimemio/_0545_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/_1105_  (.A(\soc/spimemio/_0544_ ),
    .B(\soc/spimemio/_0545_ ),
    .Y(\soc/spimemio/_0130_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/_1106_  (.A(\soc/_005_ ),
    .B(\soc/_004_ ),
    .C(\soc/_006_ ),
    .Y(\soc/spimemio/_0546_ ));
 sky130_fd_sc_hd__nand4b_1 \soc/spimemio/_1107_  (.A_N(\soc/_007_ ),
    .B(\soc/spimemio/_0546_ ),
    .C(_074_),
    .D(\soc/spimemio/config_en ),
    .Y(\soc/spimemio/_0131_ ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1108_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0014_ ),
    .Q(\soc/spimemio/buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1109_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0015_ ),
    .Q(\soc/spimemio/buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1110_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0016_ ),
    .Q(\soc/spimemio/buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1111_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0017_ ),
    .Q(\soc/spimemio/buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1112_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0018_ ),
    .Q(\soc/spimemio/buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1113_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0019_ ),
    .Q(\soc/spimemio/buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1114_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0020_ ),
    .Q(\soc/spimemio/buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1115_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0021_ ),
    .Q(\soc/spimemio/buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1116_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0022_ ),
    .Q(\soc/spimemio/din_tag[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1117_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0023_ ),
    .Q(\soc/spimemio/din_tag[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1118_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0024_ ),
    .Q(\soc/spimemio/din_tag[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1119_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0000_ ),
    .Q(\soc/spimemio/state[0] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1120_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0004_ ),
    .Q(\soc/spimemio/state[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1121_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0005_ ),
    .Q(\soc/spimemio/state[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1122_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0006_ ),
    .Q(\soc/spimemio/state[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1123_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0007_ ),
    .Q(\soc/spimemio/state[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1124_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0008_ ),
    .Q(\soc/spimemio/state[5] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1125_  (.CLK(clknet_leaf_81_clk),
    .D(net734),
    .Q(\soc/spimemio/state[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1126_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0010_ ),
    .Q(\soc/spimemio/state[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1127_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0011_ ),
    .Q(\soc/spimemio/state[8] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1128_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0012_ ),
    .Q(\soc/spimemio/state[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1129_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0001_ ),
    .Q(\soc/spimemio/state[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1130_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0002_ ),
    .Q(\soc/spimemio/state[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1131_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0003_ ),
    .Q(\soc/spimemio/state[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1132_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0025_ ),
    .Q(\soc/spimemio/rd_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1133_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0026_ ),
    .Q(\soc/spimemio/rd_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1134_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0027_ ),
    .Q(\soc/spimemio/rd_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1135_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0028_ ),
    .Q(\soc/spimemio/rd_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1136_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0029_ ),
    .Q(\soc/spimemio/rd_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1137_  (.CLK(clknet_leaf_79_clk),
    .D(net749),
    .Q(\soc/spimemio/rd_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1138_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0031_ ),
    .Q(\soc/spimemio/rd_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1139_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0032_ ),
    .Q(\soc/spimemio/rd_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1140_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0033_ ),
    .Q(\soc/spimemio/rd_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1141_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0034_ ),
    .Q(\soc/spimemio/rd_addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1142_  (.CLK(clknet_leaf_79_clk),
    .D(net716),
    .Q(\soc/spimemio/rd_addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1143_  (.CLK(clknet_leaf_79_clk),
    .D(net745),
    .Q(\soc/spimemio/rd_addr[11] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1144_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0037_ ),
    .Q(\soc/spimemio/rd_addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1145_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0038_ ),
    .Q(\soc/spimemio/rd_addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1146_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0039_ ),
    .Q(\soc/spimemio/rd_addr[14] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1147_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0040_ ),
    .Q(\soc/spimemio/rd_addr[15] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1148_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0041_ ),
    .Q(\soc/spimemio/rd_addr[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1149_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0042_ ),
    .Q(\soc/spimemio/rd_addr[17] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1150_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0043_ ),
    .Q(\soc/spimemio/rd_addr[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1151_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0044_ ),
    .Q(\soc/spimemio/rd_addr[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1152_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0045_ ),
    .Q(\soc/spimemio/rd_addr[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1153_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0046_ ),
    .Q(\soc/spimemio/rd_addr[21] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1154_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0047_ ),
    .Q(\soc/spimemio/rd_addr[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1155_  (.CLK(clknet_leaf_81_clk),
    .D(net696),
    .Q(\soc/spimemio/rd_addr[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1156_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0049_ ),
    .Q(\soc/spimemio/buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1157_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0050_ ),
    .Q(\soc/spimemio/buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1158_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0051_ ),
    .Q(\soc/spimemio/buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1159_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0052_ ),
    .Q(\soc/spimemio/buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1160_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0053_ ),
    .Q(\soc/spimemio/buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1161_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0054_ ),
    .Q(\soc/spimemio/buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1162_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0055_ ),
    .Q(\soc/spimemio/buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1163_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0056_ ),
    .Q(\soc/spimemio/buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1164_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0057_ ),
    .Q(\soc/spimem_rdata[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1165_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/_0058_ ),
    .Q(\soc/spimem_rdata[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1166_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0059_ ),
    .Q(\soc/spimem_rdata[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1167_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0060_ ),
    .Q(\soc/spimem_rdata[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1168_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0061_ ),
    .Q(\soc/spimem_rdata[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1169_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0062_ ),
    .Q(\soc/spimem_rdata[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1170_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0063_ ),
    .Q(\soc/spimem_rdata[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1171_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0064_ ),
    .Q(\soc/spimem_rdata[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1172_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0065_ ),
    .Q(\soc/spimem_rdata[8] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1173_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0066_ ),
    .Q(\soc/spimem_rdata[9] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1174_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0067_ ),
    .Q(\soc/spimem_rdata[10] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1175_  (.CLK(clknet_leaf_82_clk),
    .D(net712),
    .Q(\soc/spimem_rdata[11] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1176_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0069_ ),
    .Q(\soc/spimem_rdata[12] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1177_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0070_ ),
    .Q(\soc/spimem_rdata[13] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1178_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0071_ ),
    .Q(\soc/spimem_rdata[14] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1179_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0072_ ),
    .Q(\soc/spimem_rdata[15] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1180_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0073_ ),
    .Q(\soc/spimem_rdata[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1181_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0074_ ),
    .Q(\soc/spimem_rdata[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1182_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0075_ ),
    .Q(\soc/spimem_rdata[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1183_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0076_ ),
    .Q(\soc/spimem_rdata[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1184_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0077_ ),
    .Q(\soc/spimem_rdata[20] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1185_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0078_ ),
    .Q(\soc/spimem_rdata[21] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1186_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0079_ ),
    .Q(\soc/spimem_rdata[22] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1187_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0080_ ),
    .Q(\soc/spimem_rdata[23] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1188_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0081_ ),
    .Q(\soc/spimem_rdata[24] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1189_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0082_ ),
    .Q(\soc/spimem_rdata[25] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1190_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0083_ ),
    .Q(\soc/spimem_rdata[26] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1191_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0084_ ),
    .Q(\soc/spimem_rdata[27] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1192_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0085_ ),
    .Q(\soc/spimem_rdata[28] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1193_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0086_ ),
    .Q(\soc/spimem_rdata[29] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1194_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0087_ ),
    .Q(\soc/spimem_rdata[30] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1195_  (.CLK(clknet_leaf_84_clk),
    .D(\soc/spimemio/_0088_ ),
    .Q(\soc/spimem_rdata[31] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1196_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0089_ ),
    .Q(\soc/spimemio/xfer_resetn ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1197_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0090_ ),
    .Q(\soc/spimemio/din_valid ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1198_  (.CLK(clknet_leaf_81_clk),
    .D(net738),
    .Q(\soc/spimemio/din_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1199_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/_0092_ ),
    .Q(\soc/spimemio/din_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1200_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0093_ ),
    .Q(\soc/spimemio/din_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1201_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/_0094_ ),
    .Q(\soc/spimemio/din_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1202_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/_0095_ ),
    .Q(\soc/spimemio/din_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1203_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0096_ ),
    .Q(\soc/spimemio/din_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1204_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0097_ ),
    .Q(\soc/spimemio/din_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1205_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0098_ ),
    .Q(\soc/spimemio/din_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1206_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0099_ ),
    .Q(\soc/spimemio/din_qspi ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1207_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0100_ ),
    .Q(\soc/spimemio/din_rd ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1208_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0101_ ),
    .Q(\soc/spimemio/din_ddr ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1209_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0102_ ),
    .Q(\soc/spimemio/buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1210_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/_0103_ ),
    .Q(\soc/spimemio/buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1211_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0104_ ),
    .Q(\soc/spimemio/buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1212_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0105_ ),
    .Q(\soc/spimemio/buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1213_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0106_ ),
    .Q(\soc/spimemio/buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1214_  (.CLK(clknet_leaf_83_clk),
    .D(\soc/spimemio/_0107_ ),
    .Q(\soc/spimemio/buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1215_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0108_ ),
    .Q(\soc/spimemio/buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1216_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/_0109_ ),
    .Q(\soc/spimemio/buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1217_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/_0110_ ),
    .Q(\soc/spimemio/rd_valid ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1218_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/_0111_ ),
    .Q(\soc/spimemio/rd_wait ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1219_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0112_ ),
    .Q(\soc/spimemio/rd_inc ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1220_  (.CLK(net491),
    .D(\soc/spimemio/xfer_io0_do ),
    .Q(\soc/spimemio/xfer_io0_90 ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1221_  (.CLK(net490),
    .D(\soc/spimemio/xfer_io1_do ),
    .Q(\soc/spimemio/xfer_io1_90 ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1222_  (.CLK(net489),
    .D(\soc/spimemio/xfer_io2_do ),
    .Q(\soc/spimemio/xfer_io2_90 ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1223_  (.CLK(net488),
    .D(\soc/spimemio/xfer_io3_do ),
    .Q(\soc/spimemio/xfer_io3_90 ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1224_  (.CLK(clknet_leaf_77_clk),
    .D(\soc/spimemio/_0113_ ),
    .Q(\soc/spimemio/config_en ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1225_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/spimemio/_0114_ ),
    .Q(\soc/spimemio/config_ddr ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/_1226_  (.CLK(clknet_leaf_78_clk),
    .D(\soc/spimemio/_0115_ ),
    .Q(\soc/spimemio/config_qspi ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1227_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0116_ ),
    .Q(\soc/spimemio/config_cont ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1228_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0117_ ),
    .Q(\soc/spimemio_cfgreg_do[16] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1229_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0118_ ),
    .Q(\soc/spimemio_cfgreg_do[17] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1230_  (.CLK(clknet_leaf_79_clk),
    .D(\soc/spimemio/_0119_ ),
    .Q(\soc/spimemio_cfgreg_do[18] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1231_  (.CLK(clknet_leaf_91_clk),
    .D(\soc/spimemio/_0120_ ),
    .Q(\soc/spimemio_cfgreg_do[19] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1232_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0121_ ),
    .Q(\soc/spimemio/config_oe[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1233_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0122_ ),
    .Q(\soc/spimemio/config_oe[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1234_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0123_ ),
    .Q(\soc/spimemio/config_oe[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1235_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0124_ ),
    .Q(\soc/spimemio/config_oe[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1236_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/_0125_ ),
    .Q(\soc/spimemio/config_csb ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1237_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/_0126_ ),
    .Q(\soc/spimemio/config_clk ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1238_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/_0127_ ),
    .Q(\soc/spimemio/config_do[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1239_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/_0128_ ),
    .Q(\soc/spimemio/config_do[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1240_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/_0129_ ),
    .Q(\soc/spimemio/config_do[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/_1241_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/_0130_ ),
    .Q(\soc/spimemio/config_do[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/_1242_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/_0131_ ),
    .Q(\soc/spimemio/softreset ));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_2903__474  (.HI(net474));
 sky130_fd_sc_hd__or2_1 \soc/spimemio/xfer/_179_  (.A(\soc/spimemio/xfer/count[0] ),
    .B(\soc/spimemio/xfer/count[1] ),
    .X(\soc/spimemio/xfer/_036_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/xfer/_180_  (.A_N(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer_clk ),
    .Y(\soc/spimemio/xfer/_037_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_181_  (.A0(\soc/spimemio/xfer/count[1] ),
    .A1(\soc/spimemio/xfer/count[0] ),
    .S(\soc/spimemio/xfer/xfer_dspi ),
    .X(\soc/spimemio/xfer/_038_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/spimemio/xfer/_182_  (.A1(\soc/spimemio/xfer/_036_ ),
    .A2(\soc/spimemio/xfer/_037_ ),
    .B1(\soc/spimemio/xfer/count[3] ),
    .C1(\soc/spimemio/xfer/_038_ ),
    .Y(\soc/spimemio/xfer/_039_ ));
 sky130_fd_sc_hd__o21ai_2 \soc/spimemio/xfer/_183_  (.A1(\soc/spimemio/xfer/xfer_ddr ),
    .A2(\soc/spimemio/xfer_clk ),
    .B1(\soc/spimemio/xfer/xfer_qspi ),
    .Y(\soc/spimemio/xfer/_040_ ));
 sky130_fd_sc_hd__nor2_2 \soc/spimemio/xfer/_184_  (.A(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer/xfer_dspi ),
    .Y(\soc/spimemio/xfer/_041_ ));
 sky130_fd_sc_hd__or4_4 \soc/spimemio/xfer/_185_  (.A(\soc/spimemio/xfer/dummy_count[0] ),
    .B(\soc/spimemio/xfer/dummy_count[1] ),
    .C(\soc/spimemio/xfer/dummy_count[3] ),
    .D(\soc/spimemio/xfer/dummy_count[2] ),
    .X(\soc/spimemio/xfer/_042_ ));
 sky130_fd_sc_hd__a221oi_4 \soc/spimemio/xfer/_187_  (.A1(\soc/spimemio/xfer/count[2] ),
    .A2(\soc/spimemio/xfer/_040_ ),
    .B1(\soc/spimemio/xfer/_041_ ),
    .B2(\soc/spimemio/xfer/xfer_ddr ),
    .C1(\soc/spimemio/xfer/_042_ ),
    .Y(\soc/spimemio/xfer/_044_ ));
 sky130_fd_sc_hd__nand4_4 \soc/spimemio/xfer/_188_  (.A(\soc/spimemio/din_valid ),
    .B(\soc/spimemio/xfer_resetn ),
    .C(\soc/spimemio/xfer/_039_ ),
    .D(\soc/spimemio/xfer/_044_ ),
    .Y(\soc/spimemio/xfer/_045_ ));
 sky130_fd_sc_hd__inv_8 \soc/spimemio/xfer/_190_  (.A(\soc/spimemio/xfer/_045_ ),
    .Y(\soc/spimemio/xfer/_047_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_192_  (.A(\soc/spimemio/xfer/_039_ ),
    .B(\soc/spimemio/xfer/_044_ ),
    .Y(\soc/spimemio/xfer/_048_ ));
 sky130_fd_sc_hd__or3_1 \soc/spimemio/xfer/_193_  (.A(\soc/spimemio/xfer/fetch ),
    .B(\soc/spimemio/xfer/xfer_ddr_q ),
    .C(\soc/spimemio/xfer/_048_ ),
    .X(\soc/spimemio/xfer/_049_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/spimemio/xfer/_194_  (.A_N(\soc/spimemio/xfer/last_fetch ),
    .B(\soc/spimemio/xfer/xfer_ddr_q ),
    .C(\soc/spimemio/xfer/fetch ),
    .Y(\soc/spimemio/xfer/_050_ ));
 sky130_fd_sc_hd__inv_2 \soc/spimemio/xfer/_195_  (.A(\soc/spimemio/xfer_resetn ),
    .Y(\soc/spimemio/xfer/_051_ ));
 sky130_fd_sc_hd__a21oi_4 \soc/spimemio/xfer/_196_  (.A1(\soc/spimemio/xfer/_049_ ),
    .A2(\soc/spimemio/xfer/_050_ ),
    .B1(\soc/spimemio/xfer/_051_ ),
    .Y(\soc/spimemio/dout_valid ));
 sky130_fd_sc_hd__nor4_4 \soc/spimemio/xfer/_199_  (.A(\soc/spimemio/xfer/dummy_count[0] ),
    .B(\soc/spimemio/xfer/dummy_count[1] ),
    .C(\soc/spimemio/xfer/dummy_count[3] ),
    .D(\soc/spimemio/xfer/dummy_count[2] ),
    .Y(\soc/spimemio/xfer/_054_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/xfer/_200_  (.A(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer/obuffer[7] ),
    .C(\soc/spimemio/xfer/_054_ ),
    .X(\soc/spimemio/xfer_io3_do ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_201_  (.A(\soc/spimemio/xfer/xfer_qspi ),
    .Y(\soc/spimemio/xfer/_055_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_202_  (.A(\soc/spimemio/xfer/_055_ ),
    .B(\soc/spimemio/xfer/xfer_rd ),
    .C(\soc/spimemio/xfer/_042_ ),
    .Y(\soc/spimemio/xfer_io2_oe ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/xfer/_203_  (.A(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer/obuffer[6] ),
    .C(\soc/spimemio/xfer/_054_ ),
    .X(\soc/spimemio/xfer_io2_do ));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/xfer/_204_  (.A_N(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer/xfer_dspi ),
    .Y(\soc/spimemio/xfer/_056_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_205_  (.A(\soc/spimemio/xfer/_042_ ),
    .B(\soc/spimemio/xfer/_056_ ),
    .Y(\soc/spimemio/xfer/_057_ ));
 sky130_fd_sc_hd__a32o_1 \soc/spimemio/xfer/_206_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/xfer/obuffer[5] ),
    .A3(\soc/spimemio/xfer/_054_ ),
    .B1(\soc/spimemio/xfer/_057_ ),
    .B2(\soc/spimemio/xfer/obuffer[7] ),
    .X(\soc/spimemio/xfer_io1_do ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_207_  (.A(\soc/spimemio/xfer/xfer_rd ),
    .B(\soc/spimemio/xfer/_042_ ),
    .C(\soc/spimemio/xfer/_041_ ),
    .Y(\soc/spimemio/xfer_io1_oe ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_209_  (.A(\soc/spimemio/xfer/xfer_ddr ),
    .B(\soc/spimemio/xfer/_041_ ),
    .Y(\soc/spimemio/xfer/_059_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_210_  (.A(\soc/spimemio/xfer/_054_ ),
    .B(\soc/spimemio/xfer/_059_ ),
    .Y(\soc/spimemio/xfer/_060_ ));
 sky130_fd_sc_hd__or3_4 \soc/spimemio/xfer/_211_  (.A(\soc/spimemio/xfer/xfer_ddr ),
    .B(\soc/spimemio/xfer/xfer_qspi ),
    .C(\soc/spimemio/xfer/xfer_dspi ),
    .X(\soc/spimemio/xfer/_061_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_213_  (.A(\soc/spimemio/xfer/obuffer[7] ),
    .B(\soc/spimemio/xfer/_061_ ),
    .Y(\soc/spimemio/xfer/_063_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/xfer/_214_  (.A1(\soc/spimemio/xfer/_055_ ),
    .A2(\soc/spimemio/xfer/obuffer[4] ),
    .B1(\soc/spimemio/xfer/obuffer[6] ),
    .B2(\soc/spimemio/xfer/_056_ ),
    .Y(\soc/spimemio/xfer/_064_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_215_  (.A(\soc/spimemio/xfer/_060_ ),
    .B(\soc/spimemio/xfer/_063_ ),
    .C(\soc/spimemio/xfer/_064_ ),
    .Y(\soc/spimemio/xfer_io0_do ));
 sky130_fd_sc_hd__nor3_4 \soc/spimemio/xfer/_216_  (.A(\soc/spimemio/xfer/xfer_ddr ),
    .B(\soc/spimemio/xfer/xfer_qspi ),
    .C(\soc/spimemio/xfer/xfer_dspi ),
    .Y(\soc/spimemio/xfer/_065_ ));
 sky130_fd_sc_hd__a21o_1 \soc/spimemio/xfer/_218_  (.A1(\soc/spimemio/xfer/_054_ ),
    .A2(\soc/spimemio/xfer/_065_ ),
    .B1(\soc/spimemio/xfer_io1_oe ),
    .X(\soc/spimemio/xfer_io0_oe ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_220_  (.A(\soc/spimemio/xfer/xfer_ddr ),
    .B(\soc/spimemio/xfer/_056_ ),
    .Y(\soc/spimemio/xfer/_068_ ));
 sky130_fd_sc_hd__nor4_4 \soc/spimemio/xfer/_221_  (.A(\soc/spimemio/xfer/count[0] ),
    .B(\soc/spimemio/xfer/count[1] ),
    .C(\soc/spimemio/xfer/count[3] ),
    .D(\soc/spimemio/xfer/count[2] ),
    .Y(\soc/spimemio/xfer/_069_ ));
 sky130_fd_sc_hd__a211o_2 \soc/spimemio/xfer/_222_  (.A1(\soc/spimemio/xfer/xfer_ddr ),
    .A2(\soc/spimemio/xfer/_041_ ),
    .B1(\soc/spimemio/xfer/_069_ ),
    .C1(\soc/spimemio/xfer/_042_ ),
    .X(\soc/spimemio/xfer/_070_ ));
 sky130_fd_sc_hd__a211oi_4 \soc/spimemio/xfer/_223_  (.A1(\soc/spimemio/xfer_clk ),
    .A2(\soc/spimemio/xfer/_068_ ),
    .B1(\soc/spimemio/xfer/_070_ ),
    .C1(\soc/spimemio/xfer/_051_ ),
    .Y(\soc/spimemio/xfer/_071_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_225_  (.A(flash_io0),
    .B(\soc/spimemio/xfer/_061_ ),
    .Y(\soc/spimemio/xfer/_073_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_226_  (.A(flash_io1),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_074_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_227_  (.A(\soc/spimemio/dout_data[0] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_075_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_228_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_073_ ),
    .A3(\soc/spimemio/xfer/_074_ ),
    .B1(\soc/spimemio/xfer/_075_ ),
    .Y(\soc/spimemio/xfer/_017_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_229_  (.A(flash_io1),
    .B(\soc/spimemio/xfer/_061_ ),
    .Y(\soc/spimemio/xfer/_076_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_230_  (.A(\soc/spimemio/dout_data[0] ),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_077_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_231_  (.A(\soc/spimemio/dout_data[1] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_078_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_232_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_076_ ),
    .A3(\soc/spimemio/xfer/_077_ ),
    .B1(\soc/spimemio/xfer/_078_ ),
    .Y(\soc/spimemio/xfer/_018_ ));
 sky130_fd_sc_hd__nor2_4 \soc/spimemio/xfer/_233_  (.A(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_079_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_235_  (.A(\soc/spimemio/dout_data[0] ),
    .B(\soc/spimemio/xfer/_079_ ),
    .Y(\soc/spimemio/xfer/_081_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_236_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(flash_io2),
    .B1(\soc/spimemio/dout_data[1] ),
    .B2(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_082_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_237_  (.A(\soc/spimemio/dout_data[2] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_083_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_238_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_081_ ),
    .A3(\soc/spimemio/xfer/_082_ ),
    .B1(\soc/spimemio/xfer/_083_ ),
    .Y(\soc/spimemio/xfer/_019_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_239_  (.A(net753),
    .B(\soc/spimemio/xfer/_079_ ),
    .Y(\soc/spimemio/xfer/_084_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_240_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(flash_io3),
    .B1(net970),
    .B2(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_085_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_241_  (.A(\soc/spimemio/dout_data[3] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_086_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_242_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_084_ ),
    .A3(\soc/spimemio/xfer/_085_ ),
    .B1(\soc/spimemio/xfer/_086_ ),
    .Y(\soc/spimemio/xfer/_020_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_243_  (.A(\soc/spimemio/dout_data[3] ),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_087_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_244_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/dout_data[0] ),
    .B1(\soc/spimemio/dout_data[2] ),
    .B2(\soc/spimemio/xfer/_079_ ),
    .Y(\soc/spimemio/xfer/_088_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_245_  (.A(\soc/spimemio/dout_data[4] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_089_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_246_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_087_ ),
    .A3(\soc/spimemio/xfer/_088_ ),
    .B1(\soc/spimemio/xfer/_089_ ),
    .Y(\soc/spimemio/xfer/_021_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_247_  (.A(net886),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_090_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_248_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/dout_data[1] ),
    .B1(\soc/spimemio/dout_data[3] ),
    .B2(\soc/spimemio/xfer/_079_ ),
    .Y(\soc/spimemio/xfer/_091_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_249_  (.A(\soc/spimemio/dout_data[5] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_092_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_250_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_090_ ),
    .A3(\soc/spimemio/xfer/_091_ ),
    .B1(\soc/spimemio/xfer/_092_ ),
    .Y(\soc/spimemio/xfer/_022_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_251_  (.A(\soc/spimemio/dout_data[5] ),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_093_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_252_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/dout_data[2] ),
    .B1(net971),
    .B2(\soc/spimemio/xfer/_079_ ),
    .Y(\soc/spimemio/xfer/_094_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_253_  (.A(\soc/spimemio/dout_data[6] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_095_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_254_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_093_ ),
    .A3(\soc/spimemio/xfer/_094_ ),
    .B1(\soc/spimemio/xfer/_095_ ),
    .Y(\soc/spimemio/xfer/_023_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_255_  (.A(\soc/spimemio/dout_data[6] ),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_096_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_256_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/dout_data[3] ),
    .B1(\soc/spimemio/dout_data[5] ),
    .B2(\soc/spimemio/xfer/_079_ ),
    .Y(\soc/spimemio/xfer/_097_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_257_  (.A(\soc/spimemio/dout_data[7] ),
    .B(\soc/spimemio/xfer/_071_ ),
    .Y(\soc/spimemio/xfer/_098_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_258_  (.A1(\soc/spimemio/xfer/_071_ ),
    .A2(\soc/spimemio/xfer/_096_ ),
    .A3(\soc/spimemio/xfer/_097_ ),
    .B1(\soc/spimemio/xfer/_098_ ),
    .Y(\soc/spimemio/xfer/_024_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_259_  (.A(\soc/spimemio/xfer/obuffer[0] ),
    .Y(\soc/spimemio/xfer/_099_ ));
 sky130_fd_sc_hd__a211o_1 \soc/spimemio/xfer/_260_  (.A1(\soc/spimemio/xfer/xfer_ddr ),
    .A2(\soc/spimemio/xfer/_056_ ),
    .B1(\soc/spimemio/xfer/_069_ ),
    .C1(\soc/spimemio/xfer_clk ),
    .X(\soc/spimemio/xfer/_100_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_261_  (.A(\soc/spimemio/xfer_resetn ),
    .B(\soc/spimemio/xfer/_100_ ),
    .Y(\soc/spimemio/xfer/_101_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_262_  (.A(\soc/spimemio/xfer/_051_ ),
    .B(\soc/spimemio/xfer/_054_ ),
    .Y(\soc/spimemio/xfer/_102_ ));
 sky130_fd_sc_hd__a41oi_4 \soc/spimemio/xfer/_263_  (.A1(\soc/spimemio/din_valid ),
    .A2(\soc/spimemio/xfer_resetn ),
    .A3(\soc/spimemio/xfer/_039_ ),
    .A4(\soc/spimemio/xfer/_044_ ),
    .B1(\soc/spimemio/xfer/_102_ ),
    .Y(\soc/spimemio/xfer/_103_ ));
 sky130_fd_sc_hd__a22oi_4 \soc/spimemio/xfer/_264_  (.A1(\soc/spimemio/xfer/_045_ ),
    .A2(\soc/spimemio/xfer/_070_ ),
    .B1(\soc/spimemio/xfer/_101_ ),
    .B2(\soc/spimemio/xfer/_103_ ),
    .Y(\soc/spimemio/xfer/_104_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_265_  (.A(\soc/spimemio/din_data[0] ),
    .B(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/xfer/_105_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_266_  (.A1(\soc/spimemio/xfer/_099_ ),
    .A2(\soc/spimemio/xfer/_104_ ),
    .B1(\soc/spimemio/xfer/_105_ ),
    .Y(\soc/spimemio/xfer/_026_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_267_  (.A(\soc/spimemio/xfer/_099_ ),
    .B(\soc/spimemio/xfer/_061_ ),
    .Y(\soc/spimemio/xfer/_106_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_268_  (.A0(\soc/spimemio/din_data[1] ),
    .A1(\soc/spimemio/xfer/_106_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .X(\soc/spimemio/xfer/_107_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_269_  (.A0(\soc/spimemio/xfer/obuffer[1] ),
    .A1(\soc/spimemio/xfer/_107_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_028_ ));
 sky130_fd_sc_hd__nand2_2 \soc/spimemio/xfer/_270_  (.A(\soc/spimemio/xfer/_055_ ),
    .B(\soc/spimemio/xfer/_061_ ),
    .Y(\soc/spimemio/xfer/_108_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_271_  (.A(\soc/spimemio/xfer/obuffer[1] ),
    .B(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_109_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_272_  (.A1(\soc/spimemio/xfer/_099_ ),
    .A2(\soc/spimemio/xfer/_108_ ),
    .B1(\soc/spimemio/xfer/_109_ ),
    .Y(\soc/spimemio/xfer/_110_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_273_  (.A0(\soc/spimemio/din_data[2] ),
    .A1(\soc/spimemio/xfer/_110_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .X(\soc/spimemio/xfer/_111_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_274_  (.A0(\soc/spimemio/xfer/obuffer[2] ),
    .A1(\soc/spimemio/xfer/_111_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_029_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_275_  (.A1(\soc/spimemio/xfer/obuffer[2] ),
    .A2(\soc/spimemio/xfer/_065_ ),
    .B1(\soc/spimemio/xfer/_079_ ),
    .B2(\soc/spimemio/xfer/obuffer[1] ),
    .X(\soc/spimemio/xfer/_112_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_276_  (.A0(\soc/spimemio/din_data[3] ),
    .A1(\soc/spimemio/xfer/_112_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .X(\soc/spimemio/xfer/_113_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_277_  (.A0(\soc/spimemio/xfer/obuffer[3] ),
    .A1(\soc/spimemio/xfer/_113_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_030_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_278_  (.A(\soc/spimemio/din_data[4] ),
    .Y(\soc/spimemio/xfer/_114_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_279_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/xfer/obuffer[0] ),
    .B1(\soc/spimemio/xfer/obuffer[3] ),
    .B2(\soc/spimemio/xfer/_065_ ),
    .X(\soc/spimemio/xfer/_115_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_280_  (.A1(\soc/spimemio/xfer/obuffer[2] ),
    .A2(\soc/spimemio/xfer/_079_ ),
    .B1(\soc/spimemio/xfer/_115_ ),
    .Y(\soc/spimemio/xfer/_116_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/spimemio/xfer/_281_  (.A0(\soc/spimemio/xfer/_114_ ),
    .A1(\soc/spimemio/xfer/_116_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .Y(\soc/spimemio/xfer/_117_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_282_  (.A0(\soc/spimemio/xfer/obuffer[4] ),
    .A1(\soc/spimemio/xfer/_117_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_031_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_283_  (.A(\soc/spimemio/din_data[5] ),
    .Y(\soc/spimemio/xfer/_118_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_284_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/xfer/obuffer[1] ),
    .B1(\soc/spimemio/xfer/obuffer[4] ),
    .B2(\soc/spimemio/xfer/_065_ ),
    .X(\soc/spimemio/xfer/_119_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_285_  (.A1(\soc/spimemio/xfer/obuffer[3] ),
    .A2(\soc/spimemio/xfer/_079_ ),
    .B1(\soc/spimemio/xfer/_119_ ),
    .Y(\soc/spimemio/xfer/_120_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/spimemio/xfer/_286_  (.A0(\soc/spimemio/xfer/_118_ ),
    .A1(\soc/spimemio/xfer/_120_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .Y(\soc/spimemio/xfer/_121_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_287_  (.A0(\soc/spimemio/xfer/obuffer[5] ),
    .A1(\soc/spimemio/xfer/_121_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_032_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_288_  (.A(\soc/spimemio/din_data[6] ),
    .Y(\soc/spimemio/xfer/_122_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_289_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/xfer/obuffer[2] ),
    .B1(\soc/spimemio/xfer/obuffer[5] ),
    .B2(\soc/spimemio/xfer/_065_ ),
    .X(\soc/spimemio/xfer/_123_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_290_  (.A1(\soc/spimemio/xfer/obuffer[4] ),
    .A2(\soc/spimemio/xfer/_079_ ),
    .B1(\soc/spimemio/xfer/_123_ ),
    .Y(\soc/spimemio/xfer/_124_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/spimemio/xfer/_291_  (.A0(\soc/spimemio/xfer/_122_ ),
    .A1(\soc/spimemio/xfer/_124_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .Y(\soc/spimemio/xfer/_125_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_292_  (.A0(\soc/spimemio/xfer/obuffer[6] ),
    .A1(\soc/spimemio/xfer/_125_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_033_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_293_  (.A(\soc/spimemio/din_data[7] ),
    .Y(\soc/spimemio/xfer/_126_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_294_  (.A1(\soc/spimemio/xfer/xfer_qspi ),
    .A2(\soc/spimemio/xfer/obuffer[3] ),
    .B1(\soc/spimemio/xfer/obuffer[6] ),
    .B2(\soc/spimemio/xfer/_065_ ),
    .X(\soc/spimemio/xfer/_127_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_295_  (.A1(\soc/spimemio/xfer/obuffer[5] ),
    .A2(\soc/spimemio/xfer/_079_ ),
    .B1(\soc/spimemio/xfer/_127_ ),
    .Y(\soc/spimemio/xfer/_128_ ));
 sky130_fd_sc_hd__mux2i_1 \soc/spimemio/xfer/_296_  (.A0(\soc/spimemio/xfer/_126_ ),
    .A1(\soc/spimemio/xfer/_128_ ),
    .S(\soc/spimemio/xfer/_045_ ),
    .Y(\soc/spimemio/xfer/_129_ ));
 sky130_fd_sc_hd__mux2_1 \soc/spimemio/xfer/_297_  (.A0(\soc/spimemio/xfer/obuffer[7] ),
    .A1(\soc/spimemio/xfer/_129_ ),
    .S(\soc/spimemio/xfer/_104_ ),
    .X(\soc/spimemio/xfer/_034_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_298_  (.A(\soc/spimemio/xfer_clk ),
    .Y(\soc/spimemio/xfer/_130_ ));
 sky130_fd_sc_hd__nand3_2 \soc/spimemio/xfer/_299_  (.A(\soc/spimemio/din_valid ),
    .B(\soc/spimemio/xfer/_039_ ),
    .C(\soc/spimemio/xfer/_044_ ),
    .Y(\soc/spimemio/xfer/_131_ ));
 sky130_fd_sc_hd__nand2_2 \soc/spimemio/xfer/_300_  (.A(\soc/spimemio/xfer_resetn ),
    .B(\soc/spimemio/xfer/_131_ ),
    .Y(\soc/spimemio/xfer/_132_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_301_  (.A(\soc/spimemio/xfer_clk ),
    .B(\soc/spimemio/xfer_csb ),
    .Y(\soc/spimemio/xfer/_133_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_302_  (.A1(\soc/spimemio/xfer/_054_ ),
    .A2(\soc/spimemio/xfer/_069_ ),
    .B1(\soc/spimemio/xfer/_133_ ),
    .Y(\soc/spimemio/xfer/_134_ ));
 sky130_fd_sc_hd__a311oi_1 \soc/spimemio/xfer/_303_  (.A1(\soc/spimemio/xfer/_130_ ),
    .A2(\soc/spimemio/xfer/_054_ ),
    .A3(\soc/spimemio/xfer/_069_ ),
    .B1(\soc/spimemio/xfer/_132_ ),
    .C1(\soc/spimemio/xfer/_134_ ),
    .Y(\soc/spimemio/xfer/_002_ ));
 sky130_fd_sc_hd__a211oi_2 \soc/spimemio/xfer/_304_  (.A1(\soc/spimemio/xfer/xfer_ddr ),
    .A2(\soc/spimemio/xfer/_041_ ),
    .B1(\soc/spimemio/xfer/_069_ ),
    .C1(\soc/spimemio/xfer/_042_ ),
    .Y(\soc/spimemio/xfer/_135_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/xfer/_305_  (.A_N(\soc/spimemio/xfer/count[1] ),
    .B(\soc/spimemio/xfer_clk ),
    .Y(\soc/spimemio/xfer/_136_ ));
 sky130_fd_sc_hd__o32ai_1 \soc/spimemio/xfer/_306_  (.A1(\soc/spimemio/xfer/_130_ ),
    .A2(\soc/spimemio/xfer/_036_ ),
    .A3(\soc/spimemio/xfer/_061_ ),
    .B1(\soc/spimemio/xfer/_136_ ),
    .B2(\soc/spimemio/xfer/_108_ ),
    .Y(\soc/spimemio/xfer/_137_ ));
 sky130_fd_sc_hd__o22ai_1 \soc/spimemio/xfer/_307_  (.A1(\soc/spimemio/xfer/count[0] ),
    .A2(\soc/spimemio/xfer/_037_ ),
    .B1(\soc/spimemio/xfer/_065_ ),
    .B2(\soc/spimemio/xfer/xfer_qspi ),
    .Y(\soc/spimemio/xfer/_138_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/spimemio/xfer/_308_  (.A1(\soc/spimemio/xfer_clk ),
    .A2(\soc/spimemio/xfer/_108_ ),
    .B1(\soc/spimemio/xfer/_135_ ),
    .C1(\soc/spimemio/xfer/_138_ ),
    .Y(\soc/spimemio/xfer/_139_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_309_  (.A1(\soc/spimemio/xfer/_135_ ),
    .A2(\soc/spimemio/xfer/_137_ ),
    .B1(\soc/spimemio/xfer/_139_ ),
    .B2(\soc/spimemio/xfer/count[1] ),
    .Y(\soc/spimemio/xfer/_140_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_310_  (.A(\soc/spimemio/xfer/_132_ ),
    .B(\soc/spimemio/xfer/_140_ ),
    .Y(\soc/spimemio/xfer/_005_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_311_  (.A(\soc/spimemio/xfer/xfer_ddr ),
    .B(\soc/spimemio/xfer_clk ),
    .Y(\soc/spimemio/xfer/_141_ ));
 sky130_fd_sc_hd__and3_1 \soc/spimemio/xfer/_312_  (.A(\soc/spimemio/xfer/xfer_qspi ),
    .B(\soc/spimemio/xfer/count[2] ),
    .C(\soc/spimemio/xfer/_141_ ),
    .X(\soc/spimemio/xfer/_142_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_313_  (.A(\soc/spimemio/xfer/count[0] ),
    .B(\soc/spimemio/xfer/count[1] ),
    .C(\soc/spimemio/xfer/count[3] ),
    .Y(\soc/spimemio/xfer/_143_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_314_  (.A(\soc/spimemio/xfer/count[2] ),
    .B(\soc/spimemio/xfer/_040_ ),
    .C(\soc/spimemio/xfer/_143_ ),
    .Y(\soc/spimemio/xfer/_144_ ));
 sky130_fd_sc_hd__or3_2 \soc/spimemio/xfer/_315_  (.A(\soc/spimemio/xfer/count[2] ),
    .B(\soc/spimemio/xfer/_143_ ),
    .C(\soc/spimemio/xfer/_136_ ),
    .X(\soc/spimemio/xfer/_145_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_316_  (.A(\soc/spimemio/xfer/count[2] ),
    .B(\soc/spimemio/xfer/_136_ ),
    .Y(\soc/spimemio/xfer/_146_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_317_  (.A1(\soc/spimemio/xfer/_145_ ),
    .A2(\soc/spimemio/xfer/_146_ ),
    .B1(\soc/spimemio/xfer/_108_ ),
    .Y(\soc/spimemio/xfer/_147_ ));
 sky130_fd_sc_hd__o31ai_1 \soc/spimemio/xfer/_318_  (.A1(\soc/spimemio/xfer/_142_ ),
    .A2(\soc/spimemio/xfer/_144_ ),
    .A3(\soc/spimemio/xfer/_147_ ),
    .B1(\soc/spimemio/xfer/_135_ ),
    .Y(\soc/spimemio/xfer/_148_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_319_  (.A(\soc/spimemio/xfer/_042_ ),
    .B(\soc/spimemio/xfer/_061_ ),
    .C(\soc/spimemio/xfer/_069_ ),
    .Y(\soc/spimemio/xfer/_149_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_320_  (.A1(\soc/spimemio/xfer/count[0] ),
    .A2(\soc/spimemio/xfer/_136_ ),
    .B1(\soc/spimemio/xfer/count[2] ),
    .Y(\soc/spimemio/xfer/_150_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_321_  (.A1(\soc/spimemio/xfer/count[0] ),
    .A2(\soc/spimemio/xfer/_145_ ),
    .B1(\soc/spimemio/xfer/_150_ ),
    .Y(\soc/spimemio/xfer/_151_ ));
 sky130_fd_sc_hd__a22oi_1 \soc/spimemio/xfer/_322_  (.A1(\soc/spimemio/xfer/count[2] ),
    .A2(\soc/spimemio/xfer/_060_ ),
    .B1(\soc/spimemio/xfer/_149_ ),
    .B2(\soc/spimemio/xfer/_151_ ),
    .Y(\soc/spimemio/xfer/_152_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_323_  (.A1(\soc/spimemio/xfer/_148_ ),
    .A2(\soc/spimemio/xfer/_152_ ),
    .B1(\soc/spimemio/xfer/_132_ ),
    .Y(\soc/spimemio/xfer/_006_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_324_  (.A(\soc/spimemio/xfer_clk ),
    .B(\soc/spimemio/xfer/_149_ ),
    .Y(\soc/spimemio/xfer/_153_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/xfer/_325_  (.A(\soc/spimemio/xfer/count[0] ),
    .B(\soc/spimemio/xfer/_153_ ),
    .X(\soc/spimemio/xfer/_154_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_326_  (.A(\soc/spimemio/xfer/_132_ ),
    .B(\soc/spimemio/xfer/_154_ ),
    .Y(\soc/spimemio/xfer/_035_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_327_  (.A1(\soc/spimemio/xfer/count[0] ),
    .A2(\soc/spimemio/xfer/_145_ ),
    .B1(\soc/spimemio/xfer/_065_ ),
    .Y(\soc/spimemio/xfer/_155_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_328_  (.A1(\soc/spimemio/xfer/count[2] ),
    .A2(\soc/spimemio/xfer/_141_ ),
    .B1(\soc/spimemio/xfer/xfer_qspi ),
    .Y(\soc/spimemio/xfer/_156_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_329_  (.A1(\soc/spimemio/xfer/_145_ ),
    .A2(\soc/spimemio/xfer/_079_ ),
    .B1(\soc/spimemio/xfer/_070_ ),
    .Y(\soc/spimemio/xfer/_157_ ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/xfer/_330_  (.A(\soc/spimemio/xfer/count[3] ),
    .Y(\soc/spimemio/xfer/_158_ ));
 sky130_fd_sc_hd__a31o_1 \soc/spimemio/xfer/_331_  (.A1(\soc/spimemio/xfer/_155_ ),
    .A2(\soc/spimemio/xfer/_156_ ),
    .A3(\soc/spimemio/xfer/_157_ ),
    .B1(\soc/spimemio/xfer/_158_ ),
    .X(\soc/spimemio/xfer/_159_ ));
 sky130_fd_sc_hd__nor2_1 \soc/spimemio/xfer/_332_  (.A(\soc/spimemio/xfer/_145_ ),
    .B(\soc/spimemio/xfer/_108_ ),
    .Y(\soc/spimemio/xfer/_160_ ));
 sky130_fd_sc_hd__o211ai_1 \soc/spimemio/xfer/_333_  (.A1(\soc/spimemio/xfer/_144_ ),
    .A2(\soc/spimemio/xfer/_160_ ),
    .B1(\soc/spimemio/xfer/_158_ ),
    .C1(\soc/spimemio/xfer/_135_ ),
    .Y(\soc/spimemio/xfer/_161_ ));
 sky130_fd_sc_hd__a31oi_1 \soc/spimemio/xfer/_334_  (.A1(\soc/spimemio/xfer/_131_ ),
    .A2(\soc/spimemio/xfer/_159_ ),
    .A3(\soc/spimemio/xfer/_161_ ),
    .B1(\soc/spimemio/xfer/_051_ ),
    .Y(\soc/spimemio/xfer/_000_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_335_  (.A(\soc/spimemio/xfer_csb ),
    .B(\soc/spimemio/xfer/_131_ ),
    .Y(\soc/spimemio/xfer/_162_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_336_  (.A(\soc/spimemio/xfer_resetn ),
    .B(\soc/spimemio/xfer/_162_ ),
    .Y(\soc/spimemio/xfer/_001_ ));
 sky130_fd_sc_hd__a31oi_4 \soc/spimemio/xfer/_337_  (.A1(\soc/spimemio/din_valid ),
    .A2(\soc/spimemio/xfer/_039_ ),
    .A3(\soc/spimemio/xfer/_044_ ),
    .B1(\soc/spimemio/xfer/_051_ ),
    .Y(\soc/spimemio/xfer/_163_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_338_  (.A1(\soc/spimemio/xfer_dspi ),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_dspi ),
    .X(\soc/spimemio/xfer/_003_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_339_  (.A1(\soc/spimemio/xfer_ddr ),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_ddr ),
    .X(\soc/spimemio/xfer/_004_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/xfer/_340_  (.A(\soc/spimemio/xfer/dummy_count[0] ),
    .B(\soc/spimemio/xfer_clk ),
    .X(\soc/spimemio/xfer/_164_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_341_  (.A(\soc/spimemio/xfer/_045_ ),
    .B(\soc/spimemio/xfer/_164_ ),
    .Y(\soc/spimemio/xfer/_165_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/xfer/_342_  (.A(\soc/spimemio/din_rd ),
    .B(\soc/spimemio/din_data[0] ),
    .C(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/xfer/_166_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_343_  (.A1(\soc/spimemio/xfer/_165_ ),
    .A2(\soc/spimemio/xfer/_166_ ),
    .B1(\soc/spimemio/xfer/_103_ ),
    .Y(\soc/spimemio/xfer/_007_ ));
 sky130_fd_sc_hd__nand2b_1 \soc/spimemio/xfer/_344_  (.A_N(\soc/spimemio/xfer/dummy_count[0] ),
    .B(\soc/spimemio/xfer_clk ),
    .Y(\soc/spimemio/xfer/_167_ ));
 sky130_fd_sc_hd__xnor2_1 \soc/spimemio/xfer/_345_  (.A(\soc/spimemio/xfer/dummy_count[1] ),
    .B(\soc/spimemio/xfer/_167_ ),
    .Y(\soc/spimemio/xfer/_168_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_346_  (.A(\soc/spimemio/xfer/_045_ ),
    .B(\soc/spimemio/xfer/_168_ ),
    .Y(\soc/spimemio/xfer/_169_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/xfer/_347_  (.A(\soc/spimemio/din_rd ),
    .B(\soc/spimemio/din_data[1] ),
    .C(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/xfer/_170_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_348_  (.A1(\soc/spimemio/xfer/_169_ ),
    .A2(\soc/spimemio/xfer/_170_ ),
    .B1(\soc/spimemio/xfer/_103_ ),
    .Y(\soc/spimemio/xfer/_008_ ));
 sky130_fd_sc_hd__nor3_1 \soc/spimemio/xfer/_349_  (.A(\soc/spimemio/xfer/dummy_count[1] ),
    .B(\soc/spimemio/xfer/dummy_count[2] ),
    .C(\soc/spimemio/xfer/_167_ ),
    .Y(\soc/spimemio/xfer/_171_ ));
 sky130_fd_sc_hd__o21a_1 \soc/spimemio/xfer/_350_  (.A1(\soc/spimemio/xfer/dummy_count[1] ),
    .A2(\soc/spimemio/xfer/_167_ ),
    .B1(\soc/spimemio/xfer/dummy_count[2] ),
    .X(\soc/spimemio/xfer/_172_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_351_  (.A1(\soc/spimemio/xfer/_171_ ),
    .A2(\soc/spimemio/xfer/_172_ ),
    .B1(\soc/spimemio/xfer/_045_ ),
    .Y(\soc/spimemio/xfer/_173_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/xfer/_352_  (.A(\soc/spimemio/din_rd ),
    .B(\soc/spimemio/din_data[2] ),
    .C(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/xfer/_174_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_353_  (.A1(\soc/spimemio/xfer/_173_ ),
    .A2(\soc/spimemio/xfer/_174_ ),
    .B1(\soc/spimemio/xfer/_103_ ),
    .Y(\soc/spimemio/xfer/_009_ ));
 sky130_fd_sc_hd__xor2_1 \soc/spimemio/xfer/_354_  (.A(\soc/spimemio/xfer/dummy_count[3] ),
    .B(\soc/spimemio/xfer/_171_ ),
    .X(\soc/spimemio/xfer/_175_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_355_  (.A(\soc/spimemio/xfer/_045_ ),
    .B(\soc/spimemio/xfer/_175_ ),
    .Y(\soc/spimemio/xfer/_176_ ));
 sky130_fd_sc_hd__nand3_1 \soc/spimemio/xfer/_356_  (.A(\soc/spimemio/din_rd ),
    .B(\soc/spimemio/din_data[3] ),
    .C(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/xfer/_177_ ));
 sky130_fd_sc_hd__a21oi_1 \soc/spimemio/xfer/_357_  (.A1(\soc/spimemio/xfer/_176_ ),
    .A2(\soc/spimemio/xfer/_177_ ),
    .B1(\soc/spimemio/xfer/_103_ ),
    .Y(\soc/spimemio/xfer/_010_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_358_  (.A(net863),
    .B(\soc/spimemio/xfer/_047_ ),
    .Y(\soc/spimemio/xfer/_178_ ));
 sky130_fd_sc_hd__o21ai_0 \soc/spimemio/xfer/_359_  (.A1(\soc/spimemio/xfer/_055_ ),
    .A2(\soc/spimemio/xfer/_132_ ),
    .B1(\soc/spimemio/xfer/_178_ ),
    .Y(\soc/spimemio/xfer/_011_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_360_  (.A1(\soc/spimemio/din_rd ),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_rd ),
    .X(\soc/spimemio/xfer/_012_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_361_  (.A1(\soc/spimemio/din_tag[0] ),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_tag[0] ),
    .X(\soc/spimemio/xfer/_013_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_362_  (.A1(\soc/spimemio/din_tag[1] ),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_tag[1] ),
    .X(\soc/spimemio/xfer/_014_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_363_  (.A1(\soc/spimemio/din_tag[2] ),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_tag[2] ),
    .X(\soc/spimemio/xfer/_015_ ));
 sky130_fd_sc_hd__a22o_1 \soc/spimemio/xfer/_364_  (.A1(net472),
    .A2(\soc/spimemio/xfer/_047_ ),
    .B1(\soc/spimemio/xfer/_163_ ),
    .B2(\soc/spimemio/xfer/xfer_tag[3] ),
    .X(\soc/spimemio/xfer/_016_ ));
 sky130_fd_sc_hd__nand2_1 \soc/spimemio/xfer/_365_  (.A(\soc/spimemio/xfer_resetn ),
    .B(\soc/spimemio/xfer/_048_ ),
    .Y(\soc/spimemio/xfer/_025_ ));
 sky130_fd_sc_hd__nand3b_1 \soc/spimemio/xfer/_366_  (.A_N(\soc/spimemio/xfer/fetch ),
    .B(\soc/spimemio/xfer_resetn ),
    .C(\soc/spimemio/xfer/xfer_ddr ),
    .Y(\soc/spimemio/xfer/_027_ ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_367_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_000_ ),
    .Q(\soc/spimemio/xfer/count[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_368_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_001_ ),
    .Q(\soc/spimemio/xfer_csb ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/xfer/_369_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_002_ ),
    .Q(\soc/spimemio/xfer_clk ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_370_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_003_ ),
    .Q(\soc/spimemio/xfer/xfer_dspi ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/xfer/_371_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_004_ ),
    .Q(\soc/spimemio/xfer/xfer_ddr ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_372_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_005_ ),
    .Q(\soc/spimemio/xfer/count[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_373_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/xfer/_006_ ),
    .Q(\soc/spimemio/xfer/count[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_374_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_007_ ),
    .Q(\soc/spimemio/xfer/dummy_count[0] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_375_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_008_ ),
    .Q(\soc/spimemio/xfer/dummy_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_376_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_009_ ),
    .Q(\soc/spimemio/xfer/dummy_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_377_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_010_ ),
    .Q(\soc/spimemio/xfer/dummy_count[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/xfer/_378_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_011_ ),
    .Q(\soc/spimemio/xfer/xfer_qspi ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_379_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_012_ ),
    .Q(\soc/spimemio/xfer/xfer_rd ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_380_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/xfer/_013_ ),
    .Q(\soc/spimemio/xfer/xfer_tag[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_381_  (.CLK(clknet_leaf_81_clk),
    .D(\soc/spimemio/xfer/_014_ ),
    .Q(\soc/spimemio/xfer/xfer_tag[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_382_  (.CLK(clknet_leaf_80_clk),
    .D(\soc/spimemio/xfer/_015_ ),
    .Q(\soc/spimemio/xfer/xfer_tag[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_383_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_016_ ),
    .Q(\soc/spimemio/xfer/xfer_tag[3] ));
 sky130_fd_sc_hd__dfxtp_4 \soc/spimemio/xfer/_384_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_017_ ),
    .Q(\soc/spimemio/dout_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_385_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_018_ ),
    .Q(\soc/spimemio/dout_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_386_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_019_ ),
    .Q(\soc/spimemio/dout_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_387_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/xfer/_020_ ),
    .Q(\soc/spimemio/dout_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_388_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_021_ ),
    .Q(\soc/spimemio/dout_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_389_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/xfer/_022_ ),
    .Q(\soc/spimemio/dout_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_390_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/xfer/_023_ ),
    .Q(\soc/spimemio/dout_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_391_  (.CLK(clknet_leaf_82_clk),
    .D(\soc/spimemio/xfer/_024_ ),
    .Q(\soc/spimemio/dout_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_392_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_025_ ),
    .Q(\soc/spimemio/xfer/fetch ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_393_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/xfer_ddr ),
    .Q(\soc/spimemio/xfer/xfer_ddr_q ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_394_  (.CLK(clknet_leaf_82_clk),
    .D(net894),
    .Q(\soc/spimemio/dout_tag[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_395_  (.CLK(clknet_leaf_82_clk),
    .D(net891),
    .Q(\soc/spimemio/dout_tag[1] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_396_  (.CLK(clknet_leaf_80_clk),
    .D(net871),
    .Q(\soc/spimemio/dout_tag[2] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_397_  (.CLK(clknet_leaf_75_clk),
    .D(net870),
    .Q(\soc/spimemio/dout_tag[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_398_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_026_ ),
    .Q(\soc/spimemio/xfer/obuffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_399_  (.CLK(clknet_leaf_75_clk),
    .D(\soc/spimemio/xfer/_027_ ),
    .Q(\soc/spimemio/xfer/last_fetch ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_400_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_028_ ),
    .Q(\soc/spimemio/xfer/obuffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_401_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_029_ ),
    .Q(\soc/spimemio/xfer/obuffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_402_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_030_ ),
    .Q(\soc/spimemio/xfer/obuffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_403_  (.CLK(clknet_leaf_73_clk),
    .D(\soc/spimemio/xfer/_031_ ),
    .Q(\soc/spimemio/xfer/obuffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_404_  (.CLK(clknet_leaf_74_clk),
    .D(\soc/spimemio/xfer/_032_ ),
    .Q(\soc/spimemio/xfer/obuffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_405_  (.CLK(clknet_leaf_73_clk),
    .D(\soc/spimemio/xfer/_033_ ),
    .Q(\soc/spimemio/xfer/obuffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 \soc/spimemio/xfer/_406_  (.CLK(clknet_leaf_73_clk),
    .D(\soc/spimemio/xfer/_034_ ),
    .Q(\soc/spimemio/xfer/obuffer[7] ));
 sky130_fd_sc_hd__dfxtp_2 \soc/spimemio/xfer/_407_  (.CLK(clknet_leaf_72_clk),
    .D(\soc/spimemio/xfer/_035_ ),
    .Q(\soc/spimemio/xfer/count[0] ));
 sky130_fd_sc_hd__nand2b_4 \wave_gen_inst/_2209_  (.A_N(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/param2[4] ),
    .Y(\wave_gen_inst/_1514_ ));
 sky130_fd_sc_hd__or4_4 \wave_gen_inst/_2220_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/param2[7] ),
    .C(\wave_gen_inst/param2[8] ),
    .D(\wave_gen_inst/param2[9] ),
    .X(\wave_gen_inst/_1525_ ));
 sky130_fd_sc_hd__nor3_4 \wave_gen_inst/_2221_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/param2[11] ),
    .C(\wave_gen_inst/_1525_ ),
    .Y(\wave_gen_inst/_1526_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2223_  (.A(\wave_gen_inst/counter[11] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1528_ ));
 sky130_fd_sc_hd__inv_4 \wave_gen_inst/_2226_  (.A(\wave_gen_inst/param2[0] ),
    .Y(\wave_gen_inst/_1531_ ));
 sky130_fd_sc_hd__or3_4 \wave_gen_inst/_2228_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/param2[11] ),
    .C(\wave_gen_inst/_1525_ ),
    .X(\wave_gen_inst/_1533_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_2230_  (.A(\wave_gen_inst/_1531_ ),
    .B(\wave_gen_inst/_1533_ ),
    .Y(\wave_gen_inst/_1535_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2232_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/_1535_ ),
    .Y(\wave_gen_inst/_1537_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2233_  (.A1(\wave_gen_inst/param2[0] ),
    .A2(\wave_gen_inst/_1528_ ),
    .B1(\wave_gen_inst/_1537_ ),
    .Y(\wave_gen_inst/_1538_ ));
 sky130_fd_sc_hd__nor2_8 \wave_gen_inst/_2236_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/_1533_ ),
    .Y(\wave_gen_inst/_1541_ ));
 sky130_fd_sc_hd__a22oi_2 \wave_gen_inst/_2239_  (.A1(\wave_gen_inst/counter[10] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1541_ ),
    .B2(\wave_gen_inst/counter[9] ),
    .Y(\wave_gen_inst/_1544_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2240_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1544_ ),
    .Y(\wave_gen_inst/_1545_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2241_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1538_ ),
    .B1(\wave_gen_inst/_1545_ ),
    .Y(\wave_gen_inst/_1546_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2242_  (.A(\wave_gen_inst/_1514_ ),
    .B(\wave_gen_inst/_1546_ ),
    .Y(\wave_gen_inst/_1547_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2243_  (.A(\wave_gen_inst/param2[1] ),
    .Y(\wave_gen_inst/_1548_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2245_  (.A(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_1550_ ));
 sky130_fd_sc_hd__nand2_4 \wave_gen_inst/_2246_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1551_ ));
 sky130_fd_sc_hd__inv_6 \wave_gen_inst/_2247_  (.A(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1552_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_2249_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/param2[5] ),
    .Y(\wave_gen_inst/_1554_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2250_  (.A(\wave_gen_inst/_1552_ ),
    .B(\wave_gen_inst/_1554_ ),
    .Y(\wave_gen_inst/_1555_ ));
 sky130_fd_sc_hd__nor4_2 \wave_gen_inst/_2251_  (.A(\wave_gen_inst/_1548_ ),
    .B(\wave_gen_inst/_1550_ ),
    .C(\wave_gen_inst/_1551_ ),
    .D(\wave_gen_inst/_1555_ ),
    .Y(\wave_gen_inst/_1556_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2253_  (.A(\wave_gen_inst/counter[15] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1558_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2256_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_1535_ ),
    .Y(\wave_gen_inst/_1561_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2257_  (.A1(\wave_gen_inst/param2[0] ),
    .A2(\wave_gen_inst/_1558_ ),
    .B1(\wave_gen_inst/_1561_ ),
    .Y(\wave_gen_inst/_1562_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2261_  (.A(\wave_gen_inst/counter[13] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1566_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2262_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/_1566_ ),
    .Y(\wave_gen_inst/_1567_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2263_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1567_ ),
    .Y(\wave_gen_inst/_1568_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2264_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1568_ ),
    .Y(\wave_gen_inst/_1569_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2265_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1562_ ),
    .B1(\wave_gen_inst/_1569_ ),
    .Y(\wave_gen_inst/_1570_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_8 \wave_gen_inst/_2266_  (.A(\wave_gen_inst/param2[4] ),
    .SLEEP(\wave_gen_inst/param2[5] ),
    .X(\wave_gen_inst/_1571_ ));
 sky130_fd_sc_hd__nand2_8 \wave_gen_inst/_2267_  (.A(\wave_gen_inst/_1552_ ),
    .B(\wave_gen_inst/_1571_ ),
    .Y(\wave_gen_inst/_1572_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2269_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1570_ ),
    .B1(\wave_gen_inst/_1572_ ),
    .Y(\wave_gen_inst/_1574_ ));
 sky130_fd_sc_hd__o22ai_2 \wave_gen_inst/_2270_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1547_ ),
    .B1(\wave_gen_inst/_1556_ ),
    .B2(\wave_gen_inst/_1574_ ),
    .Y(\wave_gen_inst/_1575_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2273_  (.A(\wave_gen_inst/counter[4] ),
    .Y(\wave_gen_inst/_1578_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2275_  (.A(\wave_gen_inst/counter[3] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1580_ ));
 sky130_fd_sc_hd__o31ai_2 \wave_gen_inst/_2276_  (.A1(\wave_gen_inst/_1531_ ),
    .A2(\wave_gen_inst/_1578_ ),
    .A3(\wave_gen_inst/_1533_ ),
    .B1(\wave_gen_inst/_1580_ ),
    .Y(\wave_gen_inst/_1581_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2277_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1581_ ),
    .Y(\wave_gen_inst/_1582_ ));
 sky130_fd_sc_hd__a22o_1 \wave_gen_inst/_2281_  (.A1(\wave_gen_inst/counter[2] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1541_ ),
    .B2(\wave_gen_inst/counter[1] ),
    .X(\wave_gen_inst/_1586_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2282_  (.A(\wave_gen_inst/_1548_ ),
    .B(\wave_gen_inst/_1586_ ),
    .Y(\wave_gen_inst/_1587_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2283_  (.A(\wave_gen_inst/_1582_ ),
    .B(\wave_gen_inst/_1587_ ),
    .Y(\wave_gen_inst/_1588_ ));
 sky130_fd_sc_hd__inv_4 \wave_gen_inst/_2285_  (.A(\wave_gen_inst/counter[8] ),
    .Y(\wave_gen_inst/_1590_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2287_  (.A(\wave_gen_inst/counter[7] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1592_ ));
 sky130_fd_sc_hd__o22ai_2 \wave_gen_inst/_2288_  (.A1(\wave_gen_inst/_1590_ ),
    .A2(\wave_gen_inst/_1551_ ),
    .B1(\wave_gen_inst/_1592_ ),
    .B2(\wave_gen_inst/param2[0] ),
    .Y(\wave_gen_inst/_1593_ ));
 sky130_fd_sc_hd__a22oi_2 \wave_gen_inst/_2291_  (.A1(\wave_gen_inst/counter[6] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1541_ ),
    .B2(\wave_gen_inst/counter[5] ),
    .Y(\wave_gen_inst/_1596_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2292_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1596_ ),
    .Y(\wave_gen_inst/_1597_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2293_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1593_ ),
    .B1(\wave_gen_inst/_1597_ ),
    .Y(\wave_gen_inst/_1598_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2294_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1598_ ),
    .Y(\wave_gen_inst/_1599_ ));
 sky130_fd_sc_hd__or2_2 \wave_gen_inst/_2295_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/param2[5] ),
    .X(\wave_gen_inst/_1600_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_2296_  (.A(\wave_gen_inst/_1552_ ),
    .B(\wave_gen_inst/_1600_ ),
    .Y(\wave_gen_inst/_1601_ ));
 sky130_fd_sc_hd__o211ai_2 \wave_gen_inst/_2297_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1588_ ),
    .B1(\wave_gen_inst/_1599_ ),
    .C1(\wave_gen_inst/_1601_ ),
    .Y(\wave_gen_inst/_1602_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2301_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1606_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2302_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/_1606_ ),
    .Y(\wave_gen_inst/_1607_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2303_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1607_ ),
    .Y(\wave_gen_inst/_1608_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2306_  (.A(\wave_gen_inst/counter[17] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1611_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2308_  (.A(\wave_gen_inst/counter[18] ),
    .B(\wave_gen_inst/_1535_ ),
    .Y(\wave_gen_inst/_1613_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2309_  (.A1(\wave_gen_inst/param2[0] ),
    .A2(\wave_gen_inst/_1611_ ),
    .B1(\wave_gen_inst/_1613_ ),
    .Y(\wave_gen_inst/_1614_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2310_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1614_ ),
    .Y(\wave_gen_inst/_1615_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2311_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1608_ ),
    .B1(\wave_gen_inst/_1615_ ),
    .Y(\wave_gen_inst/_1616_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2315_  (.A(\wave_gen_inst/counter[21] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1620_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2317_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/_1535_ ),
    .Y(\wave_gen_inst/_1622_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2318_  (.A1(\wave_gen_inst/param2[0] ),
    .A2(\wave_gen_inst/_1620_ ),
    .B1(\wave_gen_inst/_1622_ ),
    .Y(\wave_gen_inst/_1623_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2322_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1627_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2323_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/_1627_ ),
    .Y(\wave_gen_inst/_1628_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_2324_  (.A1(\wave_gen_inst/counter[24] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1628_ ),
    .Y(\wave_gen_inst/_1629_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2325_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1629_ ),
    .Y(\wave_gen_inst/_1630_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2326_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1623_ ),
    .B1(\wave_gen_inst/_1630_ ),
    .Y(\wave_gen_inst/_1631_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2327_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1631_ ),
    .B1(\wave_gen_inst/_1514_ ),
    .Y(\wave_gen_inst/_1632_ ));
 sky130_fd_sc_hd__o211ai_2 \wave_gen_inst/_2330_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1616_ ),
    .B1(\wave_gen_inst/_1632_ ),
    .C1(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1635_ ));
 sky130_fd_sc_hd__nand3_4 \wave_gen_inst/_2331_  (.A(\wave_gen_inst/_1575_ ),
    .B(\wave_gen_inst/_1602_ ),
    .C(\wave_gen_inst/_1635_ ),
    .Y(\wave_gen_inst/sine_phase[0] ));
 sky130_fd_sc_hd__o2bb2a_1 \wave_gen_inst/_2332_  (.A1_N(\wave_gen_inst/counter[22] ),
    .A2_N(\wave_gen_inst/_1541_ ),
    .B1(\wave_gen_inst/_1627_ ),
    .B2(\wave_gen_inst/_1531_ ),
    .X(\wave_gen_inst/_1636_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2333_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1636_ ),
    .Y(\wave_gen_inst/_1637_ ));
 sky130_fd_sc_hd__a31oi_2 \wave_gen_inst/_2334_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/counter[24] ),
    .A3(\wave_gen_inst/_1541_ ),
    .B1(\wave_gen_inst/_1637_ ),
    .Y(\wave_gen_inst/_1638_ ));
 sky130_fd_sc_hd__o2bb2a_1 \wave_gen_inst/_2335_  (.A1_N(\wave_gen_inst/counter[20] ),
    .A2_N(\wave_gen_inst/_1541_ ),
    .B1(\wave_gen_inst/_1620_ ),
    .B2(\wave_gen_inst/_1531_ ),
    .X(\wave_gen_inst/_1639_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2336_  (.A(\wave_gen_inst/counter[18] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1640_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2337_  (.A1(\wave_gen_inst/_1531_ ),
    .A2(\wave_gen_inst/_1606_ ),
    .B1(\wave_gen_inst/_1640_ ),
    .Y(\wave_gen_inst/_1641_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2338_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1641_ ),
    .Y(\wave_gen_inst/_1642_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2339_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1639_ ),
    .B1(\wave_gen_inst/_1642_ ),
    .Y(\wave_gen_inst/_1643_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2340_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1643_ ),
    .B1(\wave_gen_inst/_1571_ ),
    .Y(\wave_gen_inst/_1644_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2341_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1638_ ),
    .B1(\wave_gen_inst/_1644_ ),
    .Y(\wave_gen_inst/_1645_ ));
 sky130_fd_sc_hd__clkinv_4 \wave_gen_inst/_2342_  (.A(\wave_gen_inst/counter[9] ),
    .Y(\wave_gen_inst/_1646_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2344_  (.A(\wave_gen_inst/counter[8] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1648_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2345_  (.A1(\wave_gen_inst/_1646_ ),
    .A2(\wave_gen_inst/_1551_ ),
    .B1(\wave_gen_inst/_1648_ ),
    .Y(\wave_gen_inst/_1649_ ));
 sky130_fd_sc_hd__o2bb2a_1 \wave_gen_inst/_2346_  (.A1_N(\wave_gen_inst/counter[6] ),
    .A2_N(\wave_gen_inst/_1541_ ),
    .B1(\wave_gen_inst/_1592_ ),
    .B2(\wave_gen_inst/_1531_ ),
    .X(\wave_gen_inst/_1650_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2347_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1650_ ),
    .Y(\wave_gen_inst/_1651_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2348_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1649_ ),
    .B1(\wave_gen_inst/_1651_ ),
    .Y(\wave_gen_inst/_1652_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2349_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/_1578_ ),
    .C(\wave_gen_inst/_1533_ ),
    .Y(\wave_gen_inst/_1653_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2350_  (.A1(\wave_gen_inst/counter[5] ),
    .A2(\wave_gen_inst/_1535_ ),
    .B1(\wave_gen_inst/_1653_ ),
    .Y(\wave_gen_inst/_1654_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2351_  (.A(\wave_gen_inst/counter[3] ),
    .Y(\wave_gen_inst/_1655_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2352_  (.A(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1656_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2353_  (.A1(\wave_gen_inst/_1655_ ),
    .A2(\wave_gen_inst/_1551_ ),
    .B1(\wave_gen_inst/_1656_ ),
    .Y(\wave_gen_inst/_1657_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2354_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1657_ ),
    .Y(\wave_gen_inst/_1658_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2355_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1654_ ),
    .B1(\wave_gen_inst/_1658_ ),
    .Y(\wave_gen_inst/_1659_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2356_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1659_ ),
    .Y(\wave_gen_inst/_1660_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_2357_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1652_ ),
    .B1(\wave_gen_inst/_1660_ ),
    .C1(\wave_gen_inst/_1600_ ),
    .Y(\wave_gen_inst/_1661_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2358_  (.A1(\wave_gen_inst/_1645_ ),
    .A2(\wave_gen_inst/_1661_ ),
    .B1(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1662_ ));
 sky130_fd_sc_hd__inv_6 \wave_gen_inst/_2359_  (.A(\wave_gen_inst/param2[2] ),
    .Y(\wave_gen_inst/_1663_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2361_  (.A(\wave_gen_inst/counter[14] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1665_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2362_  (.A1(\wave_gen_inst/_1531_ ),
    .A2(\wave_gen_inst/_1558_ ),
    .B1(\wave_gen_inst/_1665_ ),
    .Y(\wave_gen_inst/_1666_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2363_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1667_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2364_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/counter[17] ),
    .C(\wave_gen_inst/_1526_ ),
    .Y(\wave_gen_inst/_1668_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2365_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1667_ ),
    .C(\wave_gen_inst/_1668_ ),
    .Y(\wave_gen_inst/_1669_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2366_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1666_ ),
    .B1(\wave_gen_inst/_1669_ ),
    .Y(\wave_gen_inst/_1670_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2367_  (.A(\wave_gen_inst/counter[1] ),
    .Y(\wave_gen_inst/_1671_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2368_  (.A(\wave_gen_inst/_1531_ ),
    .B(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_1672_ ));
 sky130_fd_sc_hd__o22ai_2 \wave_gen_inst/_2369_  (.A1(\wave_gen_inst/_1671_ ),
    .A2(\wave_gen_inst/_1551_ ),
    .B1(\wave_gen_inst/_1672_ ),
    .B2(\wave_gen_inst/_1533_ ),
    .Y(\wave_gen_inst/_1673_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2370_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1554_ ),
    .C(\wave_gen_inst/_1673_ ),
    .Y(\wave_gen_inst/_1674_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2371_  (.A1(\wave_gen_inst/_1514_ ),
    .A2(\wave_gen_inst/_1670_ ),
    .B1(\wave_gen_inst/_1674_ ),
    .Y(\wave_gen_inst/_1675_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2372_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1676_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2373_  (.A1(\wave_gen_inst/_1531_ ),
    .A2(\wave_gen_inst/_1566_ ),
    .B1(\wave_gen_inst/_1676_ ),
    .Y(\wave_gen_inst/_1677_ ));
 sky130_fd_sc_hd__o2bb2a_1 \wave_gen_inst/_2374_  (.A1_N(\wave_gen_inst/counter[10] ),
    .A2_N(\wave_gen_inst/_1541_ ),
    .B1(\wave_gen_inst/_1528_ ),
    .B2(\wave_gen_inst/_1531_ ),
    .X(\wave_gen_inst/_1678_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2375_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1678_ ),
    .Y(\wave_gen_inst/_1679_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2376_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1677_ ),
    .B1(\wave_gen_inst/_1679_ ),
    .Y(\wave_gen_inst/_1680_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2377_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1552_ ),
    .Y(\wave_gen_inst/_1681_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2378_  (.A1(\wave_gen_inst/_1572_ ),
    .A2(\wave_gen_inst/_1680_ ),
    .B1(\wave_gen_inst/_1681_ ),
    .Y(\wave_gen_inst/_1682_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2379_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/_1675_ ),
    .B1(\wave_gen_inst/_1682_ ),
    .Y(\wave_gen_inst/_1683_ ));
 sky130_fd_sc_hd__nand2_8 \wave_gen_inst/_2380_  (.A(\wave_gen_inst/_1662_ ),
    .B(\wave_gen_inst/_1683_ ),
    .Y(\wave_gen_inst/sine_phase[1] ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2381_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1629_ ),
    .B1(\wave_gen_inst/param2[2] ),
    .Y(\wave_gen_inst/_1684_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2382_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1608_ ),
    .Y(\wave_gen_inst/_1685_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_2383_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1623_ ),
    .B1(\wave_gen_inst/_1685_ ),
    .Y(\wave_gen_inst/_1686_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2384_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/_1686_ ),
    .B1(\wave_gen_inst/_1514_ ),
    .Y(\wave_gen_inst/_1687_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2385_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1593_ ),
    .Y(\wave_gen_inst/_1688_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2386_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1544_ ),
    .B1(\wave_gen_inst/_1688_ ),
    .Y(\wave_gen_inst/_1689_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2387_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1596_ ),
    .Y(\wave_gen_inst/_1690_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2388_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1581_ ),
    .B1(\wave_gen_inst/_1690_ ),
    .Y(\wave_gen_inst/_1691_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2389_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1691_ ),
    .Y(\wave_gen_inst/_1692_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2390_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1689_ ),
    .B1(\wave_gen_inst/_1692_ ),
    .Y(\wave_gen_inst/_1693_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \wave_gen_inst/_2391_  (.A1_N(\wave_gen_inst/_1684_ ),
    .A2_N(\wave_gen_inst/_1687_ ),
    .B1(\wave_gen_inst/_1600_ ),
    .B2(\wave_gen_inst/_1693_ ),
    .Y(\wave_gen_inst/_1694_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2392_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1568_ ),
    .Y(\wave_gen_inst/_1695_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2393_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1538_ ),
    .B1(\wave_gen_inst/_1695_ ),
    .Y(\wave_gen_inst/_1696_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2394_  (.A1(\wave_gen_inst/_1572_ ),
    .A2(\wave_gen_inst/_1696_ ),
    .B1(\wave_gen_inst/_1681_ ),
    .Y(\wave_gen_inst/_1697_ ));
 sky130_fd_sc_hd__mux2i_4 \wave_gen_inst/_2395_  (.A0(\wave_gen_inst/_1562_ ),
    .A1(\wave_gen_inst/_1614_ ),
    .S(\wave_gen_inst/param2[1] ),
    .Y(\wave_gen_inst/_1698_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_2396_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1551_ ),
    .Y(\wave_gen_inst/_1699_ ));
 sky130_fd_sc_hd__a22oi_2 \wave_gen_inst/_2397_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1586_ ),
    .B1(\wave_gen_inst/_1699_ ),
    .B2(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_1700_ ));
 sky130_fd_sc_hd__o221ai_2 \wave_gen_inst/_2398_  (.A1(\wave_gen_inst/_1514_ ),
    .A2(\wave_gen_inst/_1698_ ),
    .B1(\wave_gen_inst/_1700_ ),
    .B2(\wave_gen_inst/_1600_ ),
    .C1(\wave_gen_inst/param2[2] ),
    .Y(\wave_gen_inst/_1701_ ));
 sky130_fd_sc_hd__a22o_4 \wave_gen_inst/_2399_  (.A1(\wave_gen_inst/param2[3] ),
    .A2(\wave_gen_inst/_1694_ ),
    .B1(\wave_gen_inst/_1697_ ),
    .B2(\wave_gen_inst/_1701_ ),
    .X(\wave_gen_inst/sine_phase[2] ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2400_  (.A(\wave_gen_inst/_1667_ ),
    .B(\wave_gen_inst/_1668_ ),
    .Y(\wave_gen_inst/_1702_ ));
 sky130_fd_sc_hd__mux4_1 \wave_gen_inst/_2401_  (.A0(\wave_gen_inst/_1641_ ),
    .A1(\wave_gen_inst/_1666_ ),
    .A2(\wave_gen_inst/_1702_ ),
    .A3(\wave_gen_inst/_1677_ ),
    .S0(\wave_gen_inst/_1663_ ),
    .S1(\wave_gen_inst/_1548_ ),
    .X(\wave_gen_inst/_1703_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2402_  (.A0(\wave_gen_inst/_1639_ ),
    .A1(\wave_gen_inst/_1636_ ),
    .S(\wave_gen_inst/param2[1] ),
    .X(\wave_gen_inst/_1704_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_2403_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/param2[1] ),
    .Y(\wave_gen_inst/_1705_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_2404_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/counter[24] ),
    .C(\wave_gen_inst/_1526_ ),
    .D(\wave_gen_inst/_1705_ ),
    .Y(\wave_gen_inst/_1706_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2405_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1704_ ),
    .B1(\wave_gen_inst/_1706_ ),
    .Y(\wave_gen_inst/_1707_ ));
 sky130_fd_sc_hd__mux2i_4 \wave_gen_inst/_2406_  (.A0(\wave_gen_inst/_1703_ ),
    .A1(\wave_gen_inst/_1707_ ),
    .S(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1708_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2407_  (.A(\wave_gen_inst/_1548_ ),
    .B(\wave_gen_inst/_1654_ ),
    .Y(\wave_gen_inst/_1709_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2408_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1650_ ),
    .Y(\wave_gen_inst/_1710_ ));
 sky130_fd_sc_hd__a31oi_2 \wave_gen_inst/_2409_  (.A1(\wave_gen_inst/param2[3] ),
    .A2(\wave_gen_inst/_1709_ ),
    .A3(\wave_gen_inst/_1710_ ),
    .B1(\wave_gen_inst/param2[2] ),
    .Y(\wave_gen_inst/_1711_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_2410_  (.A1(\wave_gen_inst/_1548_ ),
    .A2(\wave_gen_inst/_1657_ ),
    .B1(\wave_gen_inst/_1552_ ),
    .X(\wave_gen_inst/_1712_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2411_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1673_ ),
    .B1(\wave_gen_inst/_1712_ ),
    .Y(\wave_gen_inst/_1713_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2412_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1678_ ),
    .Y(\wave_gen_inst/_1714_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_2413_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1649_ ),
    .B1(\wave_gen_inst/_1714_ ),
    .C1(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1715_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2414_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1713_ ),
    .C(\wave_gen_inst/_1715_ ),
    .Y(\wave_gen_inst/_1716_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2415_  (.A(\wave_gen_inst/_1554_ ),
    .B(\wave_gen_inst/_1716_ ),
    .Y(\wave_gen_inst/_1717_ ));
 sky130_fd_sc_hd__o22ai_4 \wave_gen_inst/_2416_  (.A1(\wave_gen_inst/_1514_ ),
    .A2(\wave_gen_inst/_1708_ ),
    .B1(\wave_gen_inst/_1711_ ),
    .B2(\wave_gen_inst/_1717_ ),
    .Y(\wave_gen_inst/sine_phase[3] ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2417_  (.A(\wave_gen_inst/_1572_ ),
    .B(\wave_gen_inst/_1570_ ),
    .Y(\wave_gen_inst/_1718_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_2418_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1556_ ),
    .C(\wave_gen_inst/_1718_ ),
    .X(\wave_gen_inst/_1719_ ));
 sky130_fd_sc_hd__nand2_4 \wave_gen_inst/_2419_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_1554_ ),
    .Y(\wave_gen_inst/_1720_ ));
 sky130_fd_sc_hd__nand2_4 \wave_gen_inst/_2420_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_1571_ ),
    .Y(\wave_gen_inst/_1721_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_2421_  (.A1(\wave_gen_inst/_1720_ ),
    .A2(\wave_gen_inst/_1598_ ),
    .B1(\wave_gen_inst/_1721_ ),
    .B2(\wave_gen_inst/_1631_ ),
    .Y(\wave_gen_inst/_1722_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_2422_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_1600_ ),
    .Y(\wave_gen_inst/_1723_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2423_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_1514_ ),
    .Y(\wave_gen_inst/_1724_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/_2424_  (.A1(\wave_gen_inst/_1723_ ),
    .A2(\wave_gen_inst/_1588_ ),
    .B1(\wave_gen_inst/_1616_ ),
    .B2(\wave_gen_inst/_1724_ ),
    .C1(\wave_gen_inst/_1663_ ),
    .Y(\wave_gen_inst/_1725_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2425_  (.A1(\wave_gen_inst/_1546_ ),
    .A2(\wave_gen_inst/_1720_ ),
    .B1(\wave_gen_inst/_1725_ ),
    .Y(\wave_gen_inst/_1726_ ));
 sky130_fd_sc_hd__o21a_4 \wave_gen_inst/_2426_  (.A1(\wave_gen_inst/_1719_ ),
    .A2(\wave_gen_inst/_1722_ ),
    .B1(\wave_gen_inst/_1726_ ),
    .X(\wave_gen_inst/sine_phase[4] ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2427_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1673_ ),
    .B1(\wave_gen_inst/param2[2] ),
    .Y(\wave_gen_inst/_1727_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2428_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/_1659_ ),
    .B1(\wave_gen_inst/_1723_ ),
    .Y(\wave_gen_inst/_1728_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2429_  (.A(\wave_gen_inst/_1663_ ),
    .B(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1729_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_2430_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/param2[3] ),
    .C(\wave_gen_inst/_1670_ ),
    .X(\wave_gen_inst/_1730_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2431_  (.A1(\wave_gen_inst/_1638_ ),
    .A2(\wave_gen_inst/_1729_ ),
    .B1(\wave_gen_inst/_1730_ ),
    .Y(\wave_gen_inst/_1731_ ));
 sky130_fd_sc_hd__a31o_1 \wave_gen_inst/_2432_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1552_ ),
    .A3(\wave_gen_inst/_1643_ ),
    .B1(\wave_gen_inst/_1731_ ),
    .X(\wave_gen_inst/_1732_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2433_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1680_ ),
    .Y(\wave_gen_inst/_1733_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2434_  (.A(\wave_gen_inst/_1601_ ),
    .B(\wave_gen_inst/_1733_ ),
    .Y(\wave_gen_inst/_1734_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2435_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/_1652_ ),
    .B1(\wave_gen_inst/_1734_ ),
    .Y(\wave_gen_inst/_1735_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2436_  (.A1(\wave_gen_inst/_1571_ ),
    .A2(\wave_gen_inst/_1732_ ),
    .B1(\wave_gen_inst/_1735_ ),
    .Y(\wave_gen_inst/_1736_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_2437_  (.A1(\wave_gen_inst/_1727_ ),
    .A2(\wave_gen_inst/_1728_ ),
    .B1(\wave_gen_inst/_1736_ ),
    .Y(\wave_gen_inst/sine_phase[5] ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2438_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1689_ ),
    .B1(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_1737_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2439_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1696_ ),
    .B1(\wave_gen_inst/_1737_ ),
    .Y(\wave_gen_inst/_1738_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2440_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1691_ ),
    .Y(\wave_gen_inst/_1739_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2441_  (.A(\wave_gen_inst/_1552_ ),
    .B(\wave_gen_inst/_1739_ ),
    .Y(\wave_gen_inst/_1740_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2442_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/_1700_ ),
    .B1(\wave_gen_inst/_1740_ ),
    .Y(\wave_gen_inst/_1741_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_2443_  (.A1(\wave_gen_inst/_1738_ ),
    .A2(\wave_gen_inst/_1741_ ),
    .B1(\wave_gen_inst/_1554_ ),
    .Y(\wave_gen_inst/_1742_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2444_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/param2[3] ),
    .C(\wave_gen_inst/_1698_ ),
    .Y(\wave_gen_inst/_1743_ ));
 sky130_fd_sc_hd__o32ai_2 \wave_gen_inst/_2445_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1629_ ),
    .A3(\wave_gen_inst/_1729_ ),
    .B1(\wave_gen_inst/_1686_ ),
    .B2(\wave_gen_inst/_1681_ ),
    .Y(\wave_gen_inst/_1744_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2446_  (.A1(\wave_gen_inst/_1743_ ),
    .A2(\wave_gen_inst/_1744_ ),
    .B1(\wave_gen_inst/_1571_ ),
    .Y(\wave_gen_inst/_1745_ ));
 sky130_fd_sc_hd__nand2_8 \wave_gen_inst/_2447_  (.A(\wave_gen_inst/_1742_ ),
    .B(\wave_gen_inst/_1745_ ),
    .Y(\wave_gen_inst/sine_phase[6] ));
 sky130_fd_sc_hd__nor4_4 \wave_gen_inst/_2448_  (.A(net408),
    .B(net412),
    .C(net400),
    .D(net574),
    .Y(\wave_gen_inst/_1746_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2449_  (.A(net395),
    .B(\wave_gen_inst/_1746_ ),
    .Y(\wave_gen_inst/_1747_ ));
 sky130_fd_sc_hd__and2_4 \wave_gen_inst/_2450_  (.A(net388),
    .B(\wave_gen_inst/_1747_ ),
    .X(\wave_gen_inst/_1748_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \wave_gen_inst/_2454_  (.A(net12),
    .SLEEP(net11),
    .X(\wave_gen_inst/_1752_ ));
 sky130_fd_sc_hd__and2_4 \wave_gen_inst/_2455_  (.A(net13),
    .B(\wave_gen_inst/_1752_ ),
    .X(\wave_gen_inst/_1753_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2457_  (.A(net233),
    .B(\wave_gen_inst/_1753_ ),
    .Y(\wave_gen_inst/_1755_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2460_  (.A(\wave_gen_inst/sign ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1758_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2461_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1755_ ),
    .B1(\wave_gen_inst/_1758_ ),
    .Y(\wave_gen_inst/_0062_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2465_  (.A(net11),
    .B(net12),
    .Y(\wave_gen_inst/_1762_ ));
 sky130_fd_sc_hd__nor3_4 \wave_gen_inst/_2466_  (.A(net13),
    .B(\wave_gen_inst/changed ),
    .C(\wave_gen_inst/_1762_ ),
    .Y(\wave_gen_inst/_1763_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2470_  (.A(\wave_gen_inst/param2[7] ),
    .B(\wave_gen_inst/param1[7] ),
    .Y(\wave_gen_inst/_1767_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2473_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/param1[6] ),
    .Y(\wave_gen_inst/_1770_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2474_  (.A(\wave_gen_inst/_1767_ ),
    .B(\wave_gen_inst/_1770_ ),
    .Y(\wave_gen_inst/_1771_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2477_  (.A(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/param1[5] ),
    .Y(\wave_gen_inst/_1774_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2481_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/param1[4] ),
    .Y(\wave_gen_inst/_1778_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2482_  (.A(\wave_gen_inst/_1774_ ),
    .B(\wave_gen_inst/_1778_ ),
    .X(\wave_gen_inst/_1779_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2483_  (.A(\wave_gen_inst/_1771_ ),
    .B(\wave_gen_inst/_1779_ ),
    .Y(\wave_gen_inst/_1780_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2486_  (.A(\wave_gen_inst/param2[11] ),
    .B(\wave_gen_inst/param1[11] ),
    .Y(\wave_gen_inst/_1783_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2489_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/param1[10] ),
    .Y(\wave_gen_inst/_1786_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2490_  (.A(\wave_gen_inst/_1783_ ),
    .B(\wave_gen_inst/_1786_ ),
    .Y(\wave_gen_inst/_1787_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2493_  (.A(\wave_gen_inst/param2[9] ),
    .B(\wave_gen_inst/param1[9] ),
    .Y(\wave_gen_inst/_1790_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2496_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/param1[8] ),
    .Y(\wave_gen_inst/_1793_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2497_  (.A(\wave_gen_inst/_1790_ ),
    .B(\wave_gen_inst/_1793_ ),
    .X(\wave_gen_inst/_1794_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2498_  (.A(\wave_gen_inst/_1787_ ),
    .B(\wave_gen_inst/_1794_ ),
    .Y(\wave_gen_inst/_1795_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2501_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/param1[3] ),
    .Y(\wave_gen_inst/_1798_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2504_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/param1[2] ),
    .Y(\wave_gen_inst/_1801_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2505_  (.A(\wave_gen_inst/_1798_ ),
    .B(\wave_gen_inst/_1801_ ),
    .Y(\wave_gen_inst/_1802_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2508_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/param1[1] ),
    .Y(\wave_gen_inst/_1805_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2511_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/param1[0] ),
    .Y(\wave_gen_inst/_1808_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2512_  (.A(\wave_gen_inst/_1805_ ),
    .B(\wave_gen_inst/_1808_ ),
    .Y(\wave_gen_inst/_1809_ ));
 sky130_fd_sc_hd__xnor2_4 \wave_gen_inst/_2513_  (.A(\wave_gen_inst/_1802_ ),
    .B(\wave_gen_inst/_1809_ ),
    .Y(\wave_gen_inst/_1810_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2514_  (.A(\wave_gen_inst/_1795_ ),
    .B(\wave_gen_inst/_1810_ ),
    .Y(\wave_gen_inst/_1811_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2515_  (.A(\wave_gen_inst/_1780_ ),
    .B(\wave_gen_inst/_1811_ ),
    .Y(\wave_gen_inst/_1812_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2516_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/_1763_ ),
    .Y(\wave_gen_inst/_1813_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2517_  (.A1(\wave_gen_inst/_1763_ ),
    .A2(\wave_gen_inst/_1812_ ),
    .B1(\wave_gen_inst/_1813_ ),
    .Y(\wave_gen_inst/_0066_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2518_  (.A(\wave_gen_inst/param1[1] ),
    .Y(\wave_gen_inst/_1814_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2519_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/_1763_ ),
    .Y(\wave_gen_inst/_1815_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2520_  (.A1(\wave_gen_inst/_1814_ ),
    .A2(\wave_gen_inst/_1763_ ),
    .B1(\wave_gen_inst/_1815_ ),
    .Y(\wave_gen_inst/_0067_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2521_  (.A(\wave_gen_inst/param1[2] ),
    .Y(\wave_gen_inst/_1816_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2522_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/_1763_ ),
    .Y(\wave_gen_inst/_1817_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2523_  (.A1(\wave_gen_inst/_1816_ ),
    .A2(\wave_gen_inst/_1763_ ),
    .B1(\wave_gen_inst/_1817_ ),
    .Y(\wave_gen_inst/_0068_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2524_  (.A(\wave_gen_inst/param1[3] ),
    .Y(\wave_gen_inst/_1818_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2525_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/_1763_ ),
    .Y(\wave_gen_inst/_1819_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2526_  (.A1(\wave_gen_inst/_1818_ ),
    .A2(\wave_gen_inst/_1763_ ),
    .B1(\wave_gen_inst/_1819_ ),
    .Y(\wave_gen_inst/_0069_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2527_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/_1763_ ),
    .Y(\wave_gen_inst/_1820_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2528_  (.A1(\wave_gen_inst/_1818_ ),
    .A2(\wave_gen_inst/_1763_ ),
    .B1(\wave_gen_inst/_1820_ ),
    .Y(\wave_gen_inst/_0070_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2529_  (.A0(\wave_gen_inst/param1[5] ),
    .A1(net973),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0071_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2530_  (.A0(\wave_gen_inst/param1[6] ),
    .A1(\wave_gen_inst/param1[5] ),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0072_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2531_  (.A0(\wave_gen_inst/param1[7] ),
    .A1(\wave_gen_inst/param1[6] ),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0073_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2532_  (.A0(\wave_gen_inst/param1[8] ),
    .A1(\wave_gen_inst/param1[7] ),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0074_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2533_  (.A0(\wave_gen_inst/param1[9] ),
    .A1(\wave_gen_inst/param1[8] ),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0075_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2534_  (.A0(\wave_gen_inst/param1[10] ),
    .A1(\wave_gen_inst/param1[9] ),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0076_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2535_  (.A0(\wave_gen_inst/param1[11] ),
    .A1(\wave_gen_inst/param1[10] ),
    .S(\wave_gen_inst/_1763_ ),
    .X(\wave_gen_inst/_0077_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2536_  (.A(net395),
    .B(net388),
    .C(\wave_gen_inst/_1746_ ),
    .Y(\wave_gen_inst/_1821_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2537_  (.A0(net11),
    .A1(net295),
    .S(\wave_gen_inst/_1821_ ),
    .X(\wave_gen_inst/_0078_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2538_  (.A0(net12),
    .A1(net283),
    .S(\wave_gen_inst/_1821_ ),
    .X(\wave_gen_inst/_0079_ ));
 sky130_fd_sc_hd__mux2_1 \wave_gen_inst/_2539_  (.A0(net13),
    .A1(net275),
    .S(\wave_gen_inst/_1821_ ),
    .X(\wave_gen_inst/_0080_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2541_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1747_ ),
    .Y(\wave_gen_inst/_1823_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2542_  (.A(\wave_gen_inst/_1748_ ),
    .B(\wave_gen_inst/_1823_ ),
    .Y(\wave_gen_inst/_0081_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_2543_  (.A(net232),
    .B(net235),
    .C(net224),
    .D(net221),
    .X(\wave_gen_inst/_1824_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_2544_  (.A(net197),
    .B(net200),
    .C(net189),
    .D(net193),
    .Y(\wave_gen_inst/_1825_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_2545_  (.A(net210),
    .B(net213),
    .C(net204),
    .D(net207),
    .Y(\wave_gen_inst/_1826_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_2546_  (.A(net171),
    .B(net174),
    .C(net165),
    .D(net167),
    .Y(\wave_gen_inst/_1827_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_2547_  (.A(net183),
    .B(net186),
    .C(net177),
    .D(net180),
    .Y(\wave_gen_inst/_1828_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_2548_  (.A(\wave_gen_inst/_1825_ ),
    .B(\wave_gen_inst/_1826_ ),
    .C(\wave_gen_inst/_1827_ ),
    .D(\wave_gen_inst/_1828_ ),
    .Y(\wave_gen_inst/_1829_ ));
 sky130_fd_sc_hd__or4_4 \wave_gen_inst/_2549_  (.A(net228),
    .B(net217),
    .C(\wave_gen_inst/_1824_ ),
    .D(\wave_gen_inst/_1829_ ),
    .X(\wave_gen_inst/_1830_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_2550_  (.A(net263),
    .B(net241),
    .C(net249),
    .X(\wave_gen_inst/_1831_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_2551_  (.A(net253),
    .B(net260),
    .C(\wave_gen_inst/_1830_ ),
    .D(\wave_gen_inst/_1831_ ),
    .X(\wave_gen_inst/_1832_ ));
 sky130_fd_sc_hd__nand2b_4 \wave_gen_inst/_2552_  (.A_N(net13),
    .B(\wave_gen_inst/_1752_ ),
    .Y(\wave_gen_inst/_1833_ ));
 sky130_fd_sc_hd__or3_2 \wave_gen_inst/_2554_  (.A(net281),
    .B(net267),
    .C(net275),
    .X(\wave_gen_inst/_1835_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_2555_  (.A(net265),
    .B(\wave_gen_inst/_1832_ ),
    .C(\wave_gen_inst/_1833_ ),
    .D(\wave_gen_inst/_1835_ ),
    .X(\wave_gen_inst/_1836_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2556_  (.A(\wave_gen_inst/_1832_ ),
    .Y(\wave_gen_inst/_1837_ ));
 sky130_fd_sc_hd__nor3b_4 \wave_gen_inst/_2557_  (.A(net388),
    .B(\wave_gen_inst/_1746_ ),
    .C_N(net395),
    .Y(\wave_gen_inst/_1838_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2558_  (.A1(\wave_gen_inst/_1837_ ),
    .A2(\wave_gen_inst/_1833_ ),
    .B1(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1839_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2559_  (.A1(net294),
    .A2(\wave_gen_inst/_1836_ ),
    .B1(\wave_gen_inst/_1839_ ),
    .Y(\wave_gen_inst/_1840_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2561_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1842_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2562_  (.A(\wave_gen_inst/_1840_ ),
    .B(\wave_gen_inst/_1842_ ),
    .Y(\wave_gen_inst/_0082_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_2563_  (.A(net265),
    .B(\wave_gen_inst/_1832_ ),
    .C(\wave_gen_inst/_1833_ ),
    .D(\wave_gen_inst/_1835_ ),
    .Y(\wave_gen_inst/_1843_ ));
 sky130_fd_sc_hd__o32a_1 \wave_gen_inst/_2564_  (.A1(net282),
    .A2(\wave_gen_inst/_1843_ ),
    .A3(\wave_gen_inst/_1839_ ),
    .B1(\wave_gen_inst/_1838_ ),
    .B2(net821),
    .X(\wave_gen_inst/_0083_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2565_  (.A1(net849),
    .A2(\wave_gen_inst/_1838_ ),
    .B1(\wave_gen_inst/_1839_ ),
    .B2(net275),
    .X(\wave_gen_inst/_0084_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2566_  (.A1(net839),
    .A2(\wave_gen_inst/_1838_ ),
    .B1(\wave_gen_inst/_1839_ ),
    .B2(net267),
    .X(\wave_gen_inst/_0085_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2567_  (.A1(net803),
    .A2(\wave_gen_inst/_1838_ ),
    .B1(\wave_gen_inst/_1839_ ),
    .B2(net265),
    .X(\wave_gen_inst/_0086_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2569_  (.A(net263),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1845_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2570_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1846_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2571_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1845_ ),
    .B1(\wave_gen_inst/_1846_ ),
    .Y(\wave_gen_inst/_0087_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2572_  (.A(net261),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1847_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2573_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1848_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2574_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1847_ ),
    .B1(\wave_gen_inst/_1848_ ),
    .Y(\wave_gen_inst/_0088_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2575_  (.A(net253),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1849_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2576_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1850_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2577_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1849_ ),
    .B1(\wave_gen_inst/_1850_ ),
    .Y(\wave_gen_inst/_0089_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2578_  (.A(net250),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1851_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2579_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1852_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2580_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1851_ ),
    .B1(\wave_gen_inst/_1852_ ),
    .Y(\wave_gen_inst/_0090_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2581_  (.A(net242),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1853_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2582_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1854_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2583_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1853_ ),
    .B1(\wave_gen_inst/_1854_ ),
    .Y(\wave_gen_inst/_0091_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2584_  (.A(net235),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1855_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2585_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1856_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2586_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1855_ ),
    .B1(\wave_gen_inst/_1856_ ),
    .Y(\wave_gen_inst/_0092_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2587_  (.A(net233),
    .B(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_1857_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2588_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/_1838_ ),
    .Y(\wave_gen_inst/_1858_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2589_  (.A1(\wave_gen_inst/_1838_ ),
    .A2(\wave_gen_inst/_1857_ ),
    .B1(\wave_gen_inst/_1858_ ),
    .Y(\wave_gen_inst/_0093_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2590_  (.A(net239),
    .B(net247),
    .Y(\wave_gen_inst/_1859_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_2591_  (.A(net291),
    .B(net263),
    .C(net265),
    .D(\wave_gen_inst/_1835_ ),
    .X(\wave_gen_inst/_1860_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2592_  (.A(net253),
    .B(net257),
    .C(\wave_gen_inst/_1860_ ),
    .Y(\wave_gen_inst/_1861_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2593_  (.A(\wave_gen_inst/_1859_ ),
    .B(\wave_gen_inst/_1861_ ),
    .Y(\wave_gen_inst/_1862_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2594_  (.A(\wave_gen_inst/_1830_ ),
    .B(\wave_gen_inst/_1862_ ),
    .Y(\wave_gen_inst/_1863_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2595_  (.A1(net290),
    .A2(\wave_gen_inst/_1863_ ),
    .B1(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1864_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2596_  (.A1(\wave_gen_inst/_1531_ ),
    .A2(\wave_gen_inst/_1748_ ),
    .B1(\wave_gen_inst/_1864_ ),
    .Y(\wave_gen_inst/_0094_ ));
 sky130_fd_sc_hd__and3_2 \wave_gen_inst/_2597_  (.A(net13),
    .B(net233),
    .C(\wave_gen_inst/_1752_ ),
    .X(\wave_gen_inst/_1865_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2599_  (.A(net288),
    .B(\wave_gen_inst/_1865_ ),
    .Y(\wave_gen_inst/_1867_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2600_  (.A(net279),
    .B(\wave_gen_inst/_1867_ ),
    .X(\wave_gen_inst/_1868_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2601_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1869_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2602_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1868_ ),
    .B1(\wave_gen_inst/_1869_ ),
    .Y(\wave_gen_inst/_0095_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2603_  (.A1(net279),
    .A2(net287),
    .B1(\wave_gen_inst/_1865_ ),
    .Y(\wave_gen_inst/_1870_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2604_  (.A(net272),
    .B(\wave_gen_inst/_1870_ ),
    .X(\wave_gen_inst/_1871_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2605_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1872_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2606_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1871_ ),
    .B1(\wave_gen_inst/_1872_ ),
    .Y(\wave_gen_inst/_0096_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_2607_  (.A1(net280),
    .A2(net289),
    .A3(net273),
    .B1(\wave_gen_inst/_1865_ ),
    .Y(\wave_gen_inst/_1873_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2608_  (.A(net267),
    .B(\wave_gen_inst/_1873_ ),
    .X(\wave_gen_inst/_1874_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2609_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1875_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2610_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1874_ ),
    .B1(\wave_gen_inst/_1875_ ),
    .Y(\wave_gen_inst/_0097_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2611_  (.A1(net292),
    .A2(\wave_gen_inst/_1835_ ),
    .B1(\wave_gen_inst/_1865_ ),
    .Y(\wave_gen_inst/_1876_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2612_  (.A(net265),
    .B(\wave_gen_inst/_1876_ ),
    .X(\wave_gen_inst/_1877_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2613_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1878_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2614_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1877_ ),
    .B1(\wave_gen_inst/_1878_ ),
    .Y(\wave_gen_inst/_0098_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_2615_  (.A1(net293),
    .A2(net265),
    .A3(\wave_gen_inst/_1835_ ),
    .B1(\wave_gen_inst/_1865_ ),
    .Y(\wave_gen_inst/_1879_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2616_  (.A(net263),
    .B(\wave_gen_inst/_1879_ ),
    .X(\wave_gen_inst/_1880_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2617_  (.A(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1881_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2618_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1880_ ),
    .B1(\wave_gen_inst/_1881_ ),
    .Y(\wave_gen_inst/_0099_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2619_  (.A(\wave_gen_inst/_1865_ ),
    .B(\wave_gen_inst/_1860_ ),
    .Y(\wave_gen_inst/_1882_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2620_  (.A(net258),
    .B(\wave_gen_inst/_1882_ ),
    .X(\wave_gen_inst/_1883_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2621_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1884_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2622_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1883_ ),
    .B1(\wave_gen_inst/_1884_ ),
    .Y(\wave_gen_inst/_0100_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2623_  (.A1(net259),
    .A2(\wave_gen_inst/_1860_ ),
    .B1(\wave_gen_inst/_1865_ ),
    .Y(\wave_gen_inst/_1885_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2624_  (.A(net253),
    .B(\wave_gen_inst/_1885_ ),
    .X(\wave_gen_inst/_1886_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2625_  (.A(\wave_gen_inst/param2[7] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1887_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2626_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1886_ ),
    .B1(\wave_gen_inst/_1887_ ),
    .Y(\wave_gen_inst/_0101_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2627_  (.A(\wave_gen_inst/_1755_ ),
    .B(\wave_gen_inst/_1861_ ),
    .Y(\wave_gen_inst/_1888_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2628_  (.A(net246),
    .B(\wave_gen_inst/_1888_ ),
    .Y(\wave_gen_inst/_1889_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2629_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1890_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2630_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1889_ ),
    .B1(\wave_gen_inst/_1890_ ),
    .Y(\wave_gen_inst/_0102_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2631_  (.A(net248),
    .Y(\wave_gen_inst/_1891_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2632_  (.A1(\wave_gen_inst/_1891_ ),
    .A2(\wave_gen_inst/_1861_ ),
    .B1(\wave_gen_inst/_1755_ ),
    .Y(\wave_gen_inst/_1892_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2633_  (.A(net240),
    .B(\wave_gen_inst/_1892_ ),
    .Y(\wave_gen_inst/_1893_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2634_  (.A(\wave_gen_inst/param2[9] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1894_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2635_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1893_ ),
    .B1(\wave_gen_inst/_1894_ ),
    .Y(\wave_gen_inst/_0103_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2636_  (.A(\wave_gen_inst/_1865_ ),
    .B(\wave_gen_inst/_1862_ ),
    .Y(\wave_gen_inst/_1895_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2637_  (.A(net235),
    .B(\wave_gen_inst/_1895_ ),
    .X(\wave_gen_inst/_1896_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2638_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/_1748_ ),
    .Y(\wave_gen_inst/_1897_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2639_  (.A1(\wave_gen_inst/_1748_ ),
    .A2(\wave_gen_inst/_1896_ ),
    .B1(\wave_gen_inst/_1897_ ),
    .Y(\wave_gen_inst/_0104_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2640_  (.A(\wave_gen_inst/param2[11] ),
    .Y(\wave_gen_inst/_1898_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2641_  (.A1(net235),
    .A2(\wave_gen_inst/_1862_ ),
    .B1(\wave_gen_inst/_1753_ ),
    .Y(\wave_gen_inst/_1899_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2642_  (.A(net233),
    .B(\wave_gen_inst/_1748_ ),
    .C(\wave_gen_inst/_1899_ ),
    .Y(\wave_gen_inst/_1900_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2643_  (.A1(\wave_gen_inst/_1898_ ),
    .A2(\wave_gen_inst/_1748_ ),
    .B1(\wave_gen_inst/_1900_ ),
    .Y(\wave_gen_inst/_0105_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2644_  (.A(\wave_gen_inst/param1[0] ),
    .Y(\wave_gen_inst/_1901_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2645_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_1902_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2646_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_1903_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2647_  (.A(\wave_gen_inst/_1902_ ),
    .B(\wave_gen_inst/_1903_ ),
    .X(\wave_gen_inst/_1904_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2649_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_1906_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2650_  (.A(\wave_gen_inst/_1904_ ),
    .B(\wave_gen_inst/_1906_ ),
    .Y(\wave_gen_inst/_1907_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2651_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_1908_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2652_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_1909_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2654_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_1911_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2655_  (.A(\wave_gen_inst/_1908_ ),
    .B(\wave_gen_inst/_1909_ ),
    .C(\wave_gen_inst/_1911_ ),
    .X(\wave_gen_inst/_1912_ ));
 sky130_fd_sc_hd__nand4_2 \wave_gen_inst/_2658_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/param1[7] ),
    .C(\wave_gen_inst/rom_output[0] ),
    .D(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_1915_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2659_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_1916_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2660_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_1917_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2662_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_1919_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2663_  (.A(\wave_gen_inst/_1916_ ),
    .B(\wave_gen_inst/_1917_ ),
    .C(\wave_gen_inst/_1919_ ),
    .X(\wave_gen_inst/_1920_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2664_  (.A(\wave_gen_inst/_1915_ ),
    .B(\wave_gen_inst/_1920_ ),
    .X(\wave_gen_inst/_1921_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2665_  (.A(\wave_gen_inst/_1912_ ),
    .B(\wave_gen_inst/_1921_ ),
    .Y(\wave_gen_inst/_1922_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_2666_  (.A(\wave_gen_inst/_1907_ ),
    .B(\wave_gen_inst/_1922_ ),
    .X(\wave_gen_inst/_1923_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2667_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_1924_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2669_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_1926_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2670_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_1927_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2671_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_1928_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2672_  (.A(\wave_gen_inst/_1927_ ),
    .B(\wave_gen_inst/_1928_ ),
    .X(\wave_gen_inst/_1929_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2673_  (.A(\wave_gen_inst/_1926_ ),
    .B(\wave_gen_inst/_1929_ ),
    .Y(\wave_gen_inst/_1930_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2674_  (.A(\wave_gen_inst/_1924_ ),
    .B(\wave_gen_inst/_1930_ ),
    .Y(\wave_gen_inst/_1931_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2675_  (.A(\wave_gen_inst/_1916_ ),
    .B(\wave_gen_inst/_1917_ ),
    .C(\wave_gen_inst/_1919_ ),
    .X(\wave_gen_inst/_1932_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2676_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_1933_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2677_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_1934_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2679_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_1936_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2680_  (.A(\wave_gen_inst/_1933_ ),
    .B(\wave_gen_inst/_1934_ ),
    .C(\wave_gen_inst/_1936_ ),
    .X(\wave_gen_inst/_1937_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2681_  (.A(\wave_gen_inst/_1902_ ),
    .B(\wave_gen_inst/_1903_ ),
    .C(\wave_gen_inst/_1906_ ),
    .X(\wave_gen_inst/_1938_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2682_  (.A(\wave_gen_inst/_1937_ ),
    .B(\wave_gen_inst/_1938_ ),
    .Y(\wave_gen_inst/_1939_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2683_  (.A(\wave_gen_inst/_1932_ ),
    .B(\wave_gen_inst/_1939_ ),
    .X(\wave_gen_inst/_1940_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2684_  (.A(\wave_gen_inst/_1931_ ),
    .B(\wave_gen_inst/_1940_ ),
    .X(\wave_gen_inst/_1941_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2685_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_1942_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2686_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_1943_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_2688_  (.A1(\wave_gen_inst/param1[2] ),
    .A2(\wave_gen_inst/rom_output[6] ),
    .B1(\wave_gen_inst/rom_output[7] ),
    .B2(\wave_gen_inst/param1[1] ),
    .Y(\wave_gen_inst/_1945_ ));
 sky130_fd_sc_hd__o21bai_2 \wave_gen_inst/_2689_  (.A1(\wave_gen_inst/_1942_ ),
    .A2(\wave_gen_inst/_1943_ ),
    .B1_N(\wave_gen_inst/_1945_ ),
    .Y(\wave_gen_inst/_1946_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2691_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_1948_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2692_  (.A1(\wave_gen_inst/_1942_ ),
    .A2(\wave_gen_inst/_1943_ ),
    .B1(\wave_gen_inst/_1946_ ),
    .B2(\wave_gen_inst/_1948_ ),
    .X(\wave_gen_inst/_1949_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2693_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_1950_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2694_  (.A(\wave_gen_inst/_1942_ ),
    .B(\wave_gen_inst/_1950_ ),
    .Y(\wave_gen_inst/_1951_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2696_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_1953_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2697_  (.A(\wave_gen_inst/_1951_ ),
    .B(\wave_gen_inst/_1953_ ),
    .Y(\wave_gen_inst/_1954_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2698_  (.A(\wave_gen_inst/_1912_ ),
    .B(\wave_gen_inst/_1915_ ),
    .C(\wave_gen_inst/_1920_ ),
    .X(\wave_gen_inst/_1955_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2699_  (.A(\wave_gen_inst/_1954_ ),
    .B(\wave_gen_inst/_1955_ ),
    .Y(\wave_gen_inst/_1956_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2700_  (.A(\wave_gen_inst/_1949_ ),
    .B(\wave_gen_inst/_1956_ ),
    .X(\wave_gen_inst/_1957_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2701_  (.A(\wave_gen_inst/_1923_ ),
    .B(\wave_gen_inst/_1941_ ),
    .C(\wave_gen_inst/_1957_ ),
    .X(\wave_gen_inst/_1958_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_2702_  (.A(\wave_gen_inst/_1931_ ),
    .B(\wave_gen_inst/_1940_ ),
    .X(\wave_gen_inst/_1959_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_2703_  (.A(\wave_gen_inst/_1924_ ),
    .B_N(\wave_gen_inst/_1930_ ),
    .Y(\wave_gen_inst/_1960_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2704_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_1961_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2705_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_1962_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2706_  (.A(\wave_gen_inst/_1961_ ),
    .B(\wave_gen_inst/_1962_ ),
    .X(\wave_gen_inst/_1963_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2707_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_1964_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2708_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_1965_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2709_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_1966_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2710_  (.A(\wave_gen_inst/_1964_ ),
    .B(\wave_gen_inst/_1965_ ),
    .C(\wave_gen_inst/_1966_ ),
    .X(\wave_gen_inst/_1967_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2711_  (.A(\wave_gen_inst/_1963_ ),
    .B(\wave_gen_inst/_1967_ ),
    .X(\wave_gen_inst/_1968_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2712_  (.A(\wave_gen_inst/_1933_ ),
    .B(\wave_gen_inst/_1934_ ),
    .C(\wave_gen_inst/_1936_ ),
    .X(\wave_gen_inst/_1969_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2713_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_1970_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2714_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_1971_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2715_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_1972_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2716_  (.A(\wave_gen_inst/_1970_ ),
    .B(\wave_gen_inst/_1971_ ),
    .C(\wave_gen_inst/_1972_ ),
    .X(\wave_gen_inst/_1973_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2717_  (.A(\wave_gen_inst/_1927_ ),
    .B(\wave_gen_inst/_1926_ ),
    .C(\wave_gen_inst/_1928_ ),
    .X(\wave_gen_inst/_1974_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2718_  (.A(\wave_gen_inst/_1973_ ),
    .B(\wave_gen_inst/_1974_ ),
    .Y(\wave_gen_inst/_1975_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2719_  (.A(\wave_gen_inst/_1969_ ),
    .B(\wave_gen_inst/_1975_ ),
    .Y(\wave_gen_inst/_1976_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2720_  (.A(\wave_gen_inst/_1960_ ),
    .B(\wave_gen_inst/_1968_ ),
    .C(\wave_gen_inst/_1976_ ),
    .X(\wave_gen_inst/_1977_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2721_  (.A(\wave_gen_inst/_1942_ ),
    .B(\wave_gen_inst/_1950_ ),
    .C(\wave_gen_inst/_1953_ ),
    .X(\wave_gen_inst/_1978_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2722_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_1979_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2723_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_1980_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2724_  (.A(\wave_gen_inst/_1979_ ),
    .B(\wave_gen_inst/_1980_ ),
    .Y(\wave_gen_inst/_1981_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2725_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_1982_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2726_  (.A(\wave_gen_inst/_1981_ ),
    .B(\wave_gen_inst/_1982_ ),
    .Y(\wave_gen_inst/_1983_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2727_  (.A(\wave_gen_inst/_1932_ ),
    .B(\wave_gen_inst/_1937_ ),
    .C(\wave_gen_inst/_1938_ ),
    .X(\wave_gen_inst/_1984_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2728_  (.A(\wave_gen_inst/_1983_ ),
    .B(\wave_gen_inst/_1984_ ),
    .X(\wave_gen_inst/_1985_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2729_  (.A(\wave_gen_inst/_1978_ ),
    .B(\wave_gen_inst/_1985_ ),
    .Y(\wave_gen_inst/_1986_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2730_  (.A(\wave_gen_inst/_1959_ ),
    .B(\wave_gen_inst/_1977_ ),
    .C(\wave_gen_inst/_1986_ ),
    .X(\wave_gen_inst/_1987_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2731_  (.A(\wave_gen_inst/_1958_ ),
    .B(\wave_gen_inst/_1987_ ),
    .Y(\wave_gen_inst/_1988_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2732_  (.A(\wave_gen_inst/_1949_ ),
    .B(\wave_gen_inst/_1954_ ),
    .C(\wave_gen_inst/_1955_ ),
    .X(\wave_gen_inst/_1989_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2733_  (.A(\wave_gen_inst/_1958_ ),
    .B(\wave_gen_inst/_1987_ ),
    .Y(\wave_gen_inst/_1990_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_2734_  (.A1(\wave_gen_inst/_1988_ ),
    .A2(\wave_gen_inst/_1989_ ),
    .B1(\wave_gen_inst/_1990_ ),
    .X(\wave_gen_inst/_1991_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2735_  (.A(\wave_gen_inst/_1978_ ),
    .B(\wave_gen_inst/_1983_ ),
    .C(\wave_gen_inst/_1984_ ),
    .X(\wave_gen_inst/_1992_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2736_  (.A(\wave_gen_inst/_1959_ ),
    .B(\wave_gen_inst/_1977_ ),
    .C(\wave_gen_inst/_1986_ ),
    .X(\wave_gen_inst/_1993_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2737_  (.A(\wave_gen_inst/_1979_ ),
    .B(\wave_gen_inst/_1980_ ),
    .C(\wave_gen_inst/_1982_ ),
    .X(\wave_gen_inst/_1994_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2738_  (.A(\wave_gen_inst/param1[0] ),
    .B(net473),
    .Y(\wave_gen_inst/_1995_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2739_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_1996_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2740_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_1997_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2741_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_1998_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2742_  (.A(\wave_gen_inst/_1997_ ),
    .B(\wave_gen_inst/_1998_ ),
    .Y(\wave_gen_inst/_1999_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2743_  (.A1(\wave_gen_inst/_1980_ ),
    .A2(\wave_gen_inst/_1996_ ),
    .B1(\wave_gen_inst/_1999_ ),
    .Y(\wave_gen_inst/_2000_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2744_  (.A(\wave_gen_inst/_1995_ ),
    .B(\wave_gen_inst/_2000_ ),
    .Y(\wave_gen_inst/_2001_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2745_  (.A(\wave_gen_inst/_1970_ ),
    .B(\wave_gen_inst/_1971_ ),
    .Y(\wave_gen_inst/_2002_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2746_  (.A(\wave_gen_inst/_2002_ ),
    .B(\wave_gen_inst/_1972_ ),
    .Y(\wave_gen_inst/_2003_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2747_  (.A(\wave_gen_inst/_1969_ ),
    .B(\wave_gen_inst/_2003_ ),
    .C(\wave_gen_inst/_1974_ ),
    .X(\wave_gen_inst/_2004_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2748_  (.A(\wave_gen_inst/_2001_ ),
    .B(\wave_gen_inst/_2004_ ),
    .X(\wave_gen_inst/_2005_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2749_  (.A(\wave_gen_inst/_1994_ ),
    .B(\wave_gen_inst/_2005_ ),
    .Y(\wave_gen_inst/_2006_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2750_  (.A(\wave_gen_inst/_1960_ ),
    .B(\wave_gen_inst/_1968_ ),
    .C(\wave_gen_inst/_1976_ ),
    .X(\wave_gen_inst/_2007_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2751_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_2008_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2752_  (.A1(\wave_gen_inst/_1934_ ),
    .A2(\wave_gen_inst/_2008_ ),
    .B1(\wave_gen_inst/_2002_ ),
    .B2(\wave_gen_inst/_1972_ ),
    .X(\wave_gen_inst/_2009_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_2753_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .X(\wave_gen_inst/_2010_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2754_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_2011_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2755_  (.A(\wave_gen_inst/_2008_ ),
    .B(\wave_gen_inst/_2010_ ),
    .C(\wave_gen_inst/_2011_ ),
    .X(\wave_gen_inst/_2012_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2756_  (.A(\wave_gen_inst/_1964_ ),
    .B(\wave_gen_inst/_1965_ ),
    .C(\wave_gen_inst/_1966_ ),
    .X(\wave_gen_inst/_2013_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2757_  (.A(\wave_gen_inst/_2012_ ),
    .B(\wave_gen_inst/_2013_ ),
    .X(\wave_gen_inst/_2014_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2758_  (.A(\wave_gen_inst/_2009_ ),
    .B(\wave_gen_inst/_2014_ ),
    .Y(\wave_gen_inst/_2015_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2759_  (.A(\wave_gen_inst/_1963_ ),
    .B(\wave_gen_inst/_1967_ ),
    .Y(\wave_gen_inst/_2016_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2760_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2017_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2761_  (.A(\wave_gen_inst/_1924_ ),
    .B(\wave_gen_inst/_2017_ ),
    .Y(\wave_gen_inst/_2018_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2762_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_2019_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2763_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_2020_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2764_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_2021_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2765_  (.A(\wave_gen_inst/_2019_ ),
    .B(\wave_gen_inst/_2020_ ),
    .C(\wave_gen_inst/_2021_ ),
    .X(\wave_gen_inst/_2022_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2766_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_2023_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2767_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_2024_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2768_  (.A(\wave_gen_inst/_2017_ ),
    .B(\wave_gen_inst/_2023_ ),
    .C(\wave_gen_inst/_2024_ ),
    .X(\wave_gen_inst/_2025_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2769_  (.A(\wave_gen_inst/_2018_ ),
    .B(\wave_gen_inst/_2022_ ),
    .C(\wave_gen_inst/_2025_ ),
    .X(\wave_gen_inst/_2026_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2770_  (.A(\wave_gen_inst/_2016_ ),
    .B(\wave_gen_inst/_2026_ ),
    .Y(\wave_gen_inst/_2027_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2771_  (.A(\wave_gen_inst/_2015_ ),
    .B(\wave_gen_inst/_2027_ ),
    .Y(\wave_gen_inst/_2028_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2772_  (.A(\wave_gen_inst/_2007_ ),
    .B(\wave_gen_inst/_2028_ ),
    .Y(\wave_gen_inst/_2029_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2773_  (.A(\wave_gen_inst/_2006_ ),
    .B(\wave_gen_inst/_2029_ ),
    .Y(\wave_gen_inst/_2030_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2774_  (.A(\wave_gen_inst/_1992_ ),
    .B(\wave_gen_inst/_1993_ ),
    .C(\wave_gen_inst/_2030_ ),
    .X(\wave_gen_inst/_2031_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2775_  (.A(\wave_gen_inst/_1991_ ),
    .B(\wave_gen_inst/_2031_ ),
    .Y(\wave_gen_inst/_2032_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2776_  (.A(\wave_gen_inst/_2032_ ),
    .Y(\wave_gen_inst/_2033_ ));
 sky130_fd_sc_hd__a22o_1 \wave_gen_inst/_2777_  (.A1(\wave_gen_inst/param1[7] ),
    .A2(\wave_gen_inst/rom_output[0] ),
    .B1(\wave_gen_inst/rom_output[1] ),
    .B2(\wave_gen_inst/param1[6] ),
    .X(\wave_gen_inst/_2034_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2778_  (.A(\wave_gen_inst/_1915_ ),
    .B(\wave_gen_inst/_2034_ ),
    .Y(\wave_gen_inst/_2035_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2779_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_2036_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2780_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2037_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2781_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_2038_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2782_  (.A(\wave_gen_inst/_2036_ ),
    .B(\wave_gen_inst/_2037_ ),
    .C(\wave_gen_inst/_2038_ ),
    .X(\wave_gen_inst/_2039_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2783_  (.A(\wave_gen_inst/_1908_ ),
    .B(\wave_gen_inst/_1909_ ),
    .C(\wave_gen_inst/_1911_ ),
    .X(\wave_gen_inst/_2040_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2784_  (.A(\wave_gen_inst/_2039_ ),
    .B(\wave_gen_inst/_2040_ ),
    .Y(\wave_gen_inst/_2041_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_2785_  (.A(\wave_gen_inst/_2035_ ),
    .B_N(\wave_gen_inst/_2041_ ),
    .Y(\wave_gen_inst/_2042_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2786_  (.A(\wave_gen_inst/_1907_ ),
    .B(\wave_gen_inst/_1922_ ),
    .X(\wave_gen_inst/_2043_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2787_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_2044_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2788_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_2045_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2789_  (.A(\wave_gen_inst/_1943_ ),
    .B(\wave_gen_inst/_2044_ ),
    .C(\wave_gen_inst/_2045_ ),
    .X(\wave_gen_inst/_2046_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_2790_  (.A(\wave_gen_inst/_2040_ ),
    .SLEEP(\wave_gen_inst/_2039_ ),
    .X(\wave_gen_inst/_2047_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2791_  (.A(\wave_gen_inst/_1946_ ),
    .B(\wave_gen_inst/_1948_ ),
    .Y(\wave_gen_inst/_2048_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2792_  (.A(\wave_gen_inst/_2047_ ),
    .B(\wave_gen_inst/_2048_ ),
    .Y(\wave_gen_inst/_2049_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2793_  (.A(\wave_gen_inst/_2046_ ),
    .B(\wave_gen_inst/_2049_ ),
    .Y(\wave_gen_inst/_2050_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2794_  (.A(\wave_gen_inst/_2042_ ),
    .B(\wave_gen_inst/_2043_ ),
    .C(\wave_gen_inst/_2050_ ),
    .X(\wave_gen_inst/_2051_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2795_  (.A(\wave_gen_inst/_1923_ ),
    .B(\wave_gen_inst/_1941_ ),
    .C(\wave_gen_inst/_1957_ ),
    .X(\wave_gen_inst/_2052_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2796_  (.A(\wave_gen_inst/_2047_ ),
    .Y(\wave_gen_inst/_2053_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_2797_  (.A_N(\wave_gen_inst/_2046_ ),
    .B(\wave_gen_inst/_2049_ ),
    .Y(\wave_gen_inst/_2054_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2798_  (.A1(\wave_gen_inst/_2053_ ),
    .A2(\wave_gen_inst/_2048_ ),
    .B1(\wave_gen_inst/_2054_ ),
    .Y(\wave_gen_inst/_2055_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2799_  (.A(\wave_gen_inst/_2051_ ),
    .B(\wave_gen_inst/_2052_ ),
    .C(\wave_gen_inst/_2055_ ),
    .X(\wave_gen_inst/_2056_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2800_  (.A(\wave_gen_inst/_1958_ ),
    .B(\wave_gen_inst/_1987_ ),
    .C(\wave_gen_inst/_1989_ ),
    .X(\wave_gen_inst/_2057_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_2801_  (.A(\wave_gen_inst/_2056_ ),
    .B(\wave_gen_inst/_2057_ ),
    .X(\wave_gen_inst/_2058_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2802_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_2059_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2803_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2060_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2804_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_2061_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2805_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_2062_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2806_  (.A(\wave_gen_inst/_2060_ ),
    .B(\wave_gen_inst/_2061_ ),
    .C(\wave_gen_inst/_2062_ ),
    .X(\wave_gen_inst/_2063_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2807_  (.A(\wave_gen_inst/_2036_ ),
    .B(\wave_gen_inst/_2037_ ),
    .C(\wave_gen_inst/_2038_ ),
    .X(\wave_gen_inst/_2064_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2808_  (.A(\wave_gen_inst/_2063_ ),
    .B(\wave_gen_inst/_2064_ ),
    .Y(\wave_gen_inst/_2065_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2809_  (.A(\wave_gen_inst/_2059_ ),
    .B(\wave_gen_inst/_2065_ ),
    .X(\wave_gen_inst/_2066_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2810_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_2067_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2811_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_2068_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2812_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_2069_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_2813_  (.A(\wave_gen_inst/_2067_ ),
    .B(\wave_gen_inst/_2068_ ),
    .C(\wave_gen_inst/_2069_ ),
    .X(\wave_gen_inst/_2070_ ));
 sky130_fd_sc_hd__nand4_2 \wave_gen_inst/_2814_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/param1[4] ),
    .C(\wave_gen_inst/rom_output[0] ),
    .D(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2071_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2815_  (.A(\wave_gen_inst/_2060_ ),
    .B(\wave_gen_inst/_2061_ ),
    .C(\wave_gen_inst/_2062_ ),
    .X(\wave_gen_inst/_2072_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_2816_  (.A(\wave_gen_inst/_2071_ ),
    .B_N(\wave_gen_inst/_2072_ ),
    .Y(\wave_gen_inst/_2073_ ));
 sky130_fd_sc_hd__a22o_1 \wave_gen_inst/_2817_  (.A1(\wave_gen_inst/param1[2] ),
    .A2(\wave_gen_inst/rom_output[4] ),
    .B1(\wave_gen_inst/rom_output[5] ),
    .B2(\wave_gen_inst/param1[1] ),
    .X(\wave_gen_inst/_2074_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2818_  (.A1(\wave_gen_inst/_2044_ ),
    .A2(\wave_gen_inst/_2068_ ),
    .B1(\wave_gen_inst/_2074_ ),
    .Y(\wave_gen_inst/_2075_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2819_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_2076_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2820_  (.A(\wave_gen_inst/_2075_ ),
    .B(\wave_gen_inst/_2076_ ),
    .Y(\wave_gen_inst/_2077_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2821_  (.A(\wave_gen_inst/_2073_ ),
    .B(\wave_gen_inst/_2077_ ),
    .X(\wave_gen_inst/_2078_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2822_  (.A(\wave_gen_inst/_2070_ ),
    .B(\wave_gen_inst/_2078_ ),
    .Y(\wave_gen_inst/_2079_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2823_  (.A(\wave_gen_inst/_2066_ ),
    .B(\wave_gen_inst/_2079_ ),
    .Y(\wave_gen_inst/_2080_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_2824_  (.A(\wave_gen_inst/_2059_ ),
    .B_N(\wave_gen_inst/_2065_ ),
    .Y(\wave_gen_inst/_2081_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2825_  (.A(\wave_gen_inst/_2035_ ),
    .B(\wave_gen_inst/_2041_ ),
    .Y(\wave_gen_inst/_2082_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2826_  (.A(\wave_gen_inst/_2081_ ),
    .B(\wave_gen_inst/_2082_ ),
    .Y(\wave_gen_inst/_2083_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2827_  (.A1(\wave_gen_inst/_2044_ ),
    .A2(\wave_gen_inst/_2068_ ),
    .B1(\wave_gen_inst/_2075_ ),
    .B2(\wave_gen_inst/_2076_ ),
    .X(\wave_gen_inst/_2084_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_2828_  (.A(\wave_gen_inst/_2064_ ),
    .SLEEP(\wave_gen_inst/_2063_ ),
    .X(\wave_gen_inst/_2085_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2829_  (.A(\wave_gen_inst/_1943_ ),
    .B(\wave_gen_inst/_2044_ ),
    .Y(\wave_gen_inst/_2086_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2830_  (.A(\wave_gen_inst/_2086_ ),
    .B(\wave_gen_inst/_2045_ ),
    .Y(\wave_gen_inst/_2087_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2831_  (.A(\wave_gen_inst/_2085_ ),
    .B(\wave_gen_inst/_2087_ ),
    .Y(\wave_gen_inst/_2088_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2832_  (.A(\wave_gen_inst/_2084_ ),
    .B(\wave_gen_inst/_2088_ ),
    .Y(\wave_gen_inst/_2089_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2833_  (.A(\wave_gen_inst/_2083_ ),
    .B(\wave_gen_inst/_2089_ ),
    .Y(\wave_gen_inst/_2090_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2834_  (.A(\wave_gen_inst/_2073_ ),
    .Y(\wave_gen_inst/_2091_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2835_  (.A(\wave_gen_inst/_2070_ ),
    .B(\wave_gen_inst/_2091_ ),
    .C(\wave_gen_inst/_2077_ ),
    .X(\wave_gen_inst/_2092_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2836_  (.A(\wave_gen_inst/_2092_ ),
    .Y(\wave_gen_inst/_2093_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2837_  (.A(\wave_gen_inst/_2080_ ),
    .B(\wave_gen_inst/_2090_ ),
    .C(\wave_gen_inst/_2093_ ),
    .X(\wave_gen_inst/_2094_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2838_  (.A(\wave_gen_inst/_2081_ ),
    .B(\wave_gen_inst/_2082_ ),
    .C(\wave_gen_inst/_2089_ ),
    .X(\wave_gen_inst/_2095_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2839_  (.A(\wave_gen_inst/_2042_ ),
    .B(\wave_gen_inst/_2043_ ),
    .C(\wave_gen_inst/_2050_ ),
    .X(\wave_gen_inst/_2096_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2840_  (.A(\wave_gen_inst/_2085_ ),
    .Y(\wave_gen_inst/_2097_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_2841_  (.A_N(\wave_gen_inst/_2084_ ),
    .B(\wave_gen_inst/_2088_ ),
    .Y(\wave_gen_inst/_2098_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2842_  (.A1(\wave_gen_inst/_2097_ ),
    .A2(\wave_gen_inst/_2087_ ),
    .B1(\wave_gen_inst/_2098_ ),
    .Y(\wave_gen_inst/_2099_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2843_  (.A(\wave_gen_inst/_2095_ ),
    .B(\wave_gen_inst/_2096_ ),
    .C(\wave_gen_inst/_2099_ ),
    .X(\wave_gen_inst/_2100_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2844_  (.A(\wave_gen_inst/_2080_ ),
    .B(\wave_gen_inst/_2090_ ),
    .C(\wave_gen_inst/_2092_ ),
    .X(\wave_gen_inst/_2101_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2845_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_2102_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2846_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_2103_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_2847_  (.A1(\wave_gen_inst/param1[2] ),
    .A2(\wave_gen_inst/rom_output[2] ),
    .B1(\wave_gen_inst/rom_output[3] ),
    .B2(\wave_gen_inst/param1[1] ),
    .Y(\wave_gen_inst/_2104_ ));
 sky130_fd_sc_hd__o21bai_1 \wave_gen_inst/_2848_  (.A1(\wave_gen_inst/_2067_ ),
    .A2(\wave_gen_inst/_2102_ ),
    .B1_N(\wave_gen_inst/_2104_ ),
    .Y(\wave_gen_inst/_2105_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2849_  (.A1(\wave_gen_inst/_2067_ ),
    .A2(\wave_gen_inst/_2102_ ),
    .B1(\wave_gen_inst/_2103_ ),
    .B2(\wave_gen_inst/_2105_ ),
    .X(\wave_gen_inst/_2106_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2850_  (.A(\wave_gen_inst/_2067_ ),
    .B(\wave_gen_inst/_2068_ ),
    .X(\wave_gen_inst/_2107_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2851_  (.A(\wave_gen_inst/_2069_ ),
    .B(\wave_gen_inst/_2107_ ),
    .Y(\wave_gen_inst/_2108_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_2852_  (.A_N(\wave_gen_inst/_2106_ ),
    .B(\wave_gen_inst/_2108_ ),
    .Y(\wave_gen_inst/_2109_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2853_  (.A(\wave_gen_inst/_2071_ ),
    .B(\wave_gen_inst/_2072_ ),
    .Y(\wave_gen_inst/_2110_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2854_  (.A(\wave_gen_inst/_2106_ ),
    .B(\wave_gen_inst/_2108_ ),
    .Y(\wave_gen_inst/_2111_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_2855_  (.A(\wave_gen_inst/_2110_ ),
    .B(\wave_gen_inst/_2111_ ),
    .X(\wave_gen_inst/_2112_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2856_  (.A(\wave_gen_inst/_2066_ ),
    .B(\wave_gen_inst/_2070_ ),
    .C(\wave_gen_inst/_2078_ ),
    .X(\wave_gen_inst/_2113_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2857_  (.A(\wave_gen_inst/_2112_ ),
    .B(\wave_gen_inst/_2113_ ),
    .Y(\wave_gen_inst/_2114_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2858_  (.A(\wave_gen_inst/_2110_ ),
    .B(\wave_gen_inst/_2111_ ),
    .Y(\wave_gen_inst/_2115_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2859_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2116_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2860_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_2117_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2861_  (.A(\wave_gen_inst/_2102_ ),
    .B(\wave_gen_inst/_2116_ ),
    .C(\wave_gen_inst/_2117_ ),
    .X(\wave_gen_inst/_2118_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2862_  (.A(\wave_gen_inst/_2103_ ),
    .B(\wave_gen_inst/_2105_ ),
    .Y(\wave_gen_inst/_2119_ ));
 sky130_fd_sc_hd__a22o_1 \wave_gen_inst/_2863_  (.A1(\wave_gen_inst/param1[4] ),
    .A2(\wave_gen_inst/rom_output[0] ),
    .B1(\wave_gen_inst/rom_output[1] ),
    .B2(\wave_gen_inst/param1[3] ),
    .X(\wave_gen_inst/_2120_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2864_  (.A(\wave_gen_inst/_2071_ ),
    .B(\wave_gen_inst/_2120_ ),
    .Y(\wave_gen_inst/_2121_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2865_  (.A(\wave_gen_inst/_2118_ ),
    .B(\wave_gen_inst/_2119_ ),
    .C(\wave_gen_inst/_2121_ ),
    .X(\wave_gen_inst/_2122_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2866_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2123_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2867_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_2124_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2868_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_2125_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2869_  (.A(\wave_gen_inst/_2123_ ),
    .B(\wave_gen_inst/_2124_ ),
    .C(\wave_gen_inst/_2125_ ),
    .X(\wave_gen_inst/_2126_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2870_  (.A(\wave_gen_inst/_2102_ ),
    .B(\wave_gen_inst/_2116_ ),
    .C(\wave_gen_inst/_2117_ ),
    .X(\wave_gen_inst/_2127_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2871_  (.A(\wave_gen_inst/_2126_ ),
    .B(\wave_gen_inst/_2127_ ),
    .Y(\wave_gen_inst/_2128_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2872_  (.A(\wave_gen_inst/_2123_ ),
    .B(\wave_gen_inst/_2125_ ),
    .X(\wave_gen_inst/_2129_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2873_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_2130_ ));
 sky130_fd_sc_hd__a311o_1 \wave_gen_inst/_2874_  (.A1(\wave_gen_inst/param1[2] ),
    .A2(\wave_gen_inst/rom_output[0] ),
    .A3(\wave_gen_inst/_2124_ ),
    .B1(\wave_gen_inst/_2130_ ),
    .C1(\wave_gen_inst/_2123_ ),
    .X(\wave_gen_inst/_2131_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2875_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[0] ),
    .Y(\wave_gen_inst/_2132_ ));
 sky130_fd_sc_hd__a311oi_2 \wave_gen_inst/_2876_  (.A1(\wave_gen_inst/param1[0] ),
    .A2(\wave_gen_inst/rom_output[2] ),
    .A3(\wave_gen_inst/_2129_ ),
    .B1(\wave_gen_inst/_2131_ ),
    .C1(\wave_gen_inst/_2132_ ),
    .Y(\wave_gen_inst/_2133_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_2877_  (.A1(\wave_gen_inst/param1[0] ),
    .A2(\wave_gen_inst/rom_output[2] ),
    .A3(\wave_gen_inst/_2129_ ),
    .B1(\wave_gen_inst/_2131_ ),
    .Y(\wave_gen_inst/_2134_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2878_  (.A1(\wave_gen_inst/_2126_ ),
    .A2(\wave_gen_inst/_2127_ ),
    .B1(\wave_gen_inst/_2132_ ),
    .Y(\wave_gen_inst/_2135_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2879_  (.A(\wave_gen_inst/_2126_ ),
    .B(\wave_gen_inst/_2127_ ),
    .Y(\wave_gen_inst/_2136_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_2880_  (.A1(\wave_gen_inst/_2134_ ),
    .A2(\wave_gen_inst/_2135_ ),
    .B1(\wave_gen_inst/_2133_ ),
    .B2(\wave_gen_inst/_2136_ ),
    .Y(\wave_gen_inst/_2137_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2881_  (.A(\wave_gen_inst/_2118_ ),
    .B(\wave_gen_inst/_2119_ ),
    .C(\wave_gen_inst/_2121_ ),
    .X(\wave_gen_inst/_2138_ ));
 sky130_fd_sc_hd__o2bb2a_1 \wave_gen_inst/_2882_  (.A1_N(\wave_gen_inst/_2128_ ),
    .A2_N(\wave_gen_inst/_2133_ ),
    .B1(\wave_gen_inst/_2137_ ),
    .B2(\wave_gen_inst/_2138_ ),
    .X(\wave_gen_inst/_2139_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2883_  (.A(\wave_gen_inst/_2115_ ),
    .B(\wave_gen_inst/_2122_ ),
    .C(\wave_gen_inst/_2139_ ),
    .X(\wave_gen_inst/_2140_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2884_  (.A(\wave_gen_inst/_2109_ ),
    .B(\wave_gen_inst/_2114_ ),
    .C(\wave_gen_inst/_2140_ ),
    .Y(\wave_gen_inst/_2141_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2885_  (.A(\wave_gen_inst/_2112_ ),
    .B(\wave_gen_inst/_2113_ ),
    .Y(\wave_gen_inst/_2142_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2886_  (.A1(\wave_gen_inst/_2109_ ),
    .A2(\wave_gen_inst/_2140_ ),
    .B1(\wave_gen_inst/_2142_ ),
    .Y(\wave_gen_inst/_2143_ ));
 sky130_fd_sc_hd__o2111ai_2 \wave_gen_inst/_2887_  (.A1(\wave_gen_inst/_2094_ ),
    .A2(\wave_gen_inst/_2100_ ),
    .B1(\wave_gen_inst/_2101_ ),
    .C1(\wave_gen_inst/_2141_ ),
    .D1(\wave_gen_inst/_2143_ ),
    .Y(\wave_gen_inst/_2144_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2888_  (.A(\wave_gen_inst/_2095_ ),
    .B(\wave_gen_inst/_2096_ ),
    .C(\wave_gen_inst/_2099_ ),
    .X(\wave_gen_inst/_2145_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_2889_  (.A(\wave_gen_inst/_2051_ ),
    .B(\wave_gen_inst/_2052_ ),
    .C(\wave_gen_inst/_2055_ ),
    .X(\wave_gen_inst/_2146_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_2890_  (.A1(\wave_gen_inst/_2094_ ),
    .A2(\wave_gen_inst/_2100_ ),
    .B1(\wave_gen_inst/_2145_ ),
    .B2(\wave_gen_inst/_2146_ ),
    .Y(\wave_gen_inst/_2147_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_2891_  (.A1(\wave_gen_inst/_2056_ ),
    .A2(\wave_gen_inst/_2057_ ),
    .B1(\wave_gen_inst/_2145_ ),
    .B2(\wave_gen_inst/_2146_ ),
    .Y(\wave_gen_inst/_2148_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_2892_  (.A1(\wave_gen_inst/_2144_ ),
    .A2(\wave_gen_inst/_2147_ ),
    .B1(\wave_gen_inst/_2148_ ),
    .Y(\wave_gen_inst/_2149_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2893_  (.A(\wave_gen_inst/_1991_ ),
    .B(\wave_gen_inst/_2031_ ),
    .X(\wave_gen_inst/_2150_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_2894_  (.A1(\wave_gen_inst/_2058_ ),
    .A2(\wave_gen_inst/_2149_ ),
    .B1(\wave_gen_inst/_2150_ ),
    .Y(\wave_gen_inst/_2151_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2895_  (.A(\wave_gen_inst/_2033_ ),
    .B(\wave_gen_inst/_2151_ ),
    .Y(\wave_gen_inst/_2152_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2896_  (.A(\wave_gen_inst/_1993_ ),
    .Y(\wave_gen_inst/_2153_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_2897_  (.A(\wave_gen_inst/_1992_ ),
    .B(\wave_gen_inst/_2153_ ),
    .C(\wave_gen_inst/_2030_ ),
    .X(\wave_gen_inst/_2154_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2898_  (.A(\wave_gen_inst/_1994_ ),
    .B(\wave_gen_inst/_2001_ ),
    .C(\wave_gen_inst/_2004_ ),
    .X(\wave_gen_inst/_2155_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2899_  (.A(\wave_gen_inst/_2028_ ),
    .Y(\wave_gen_inst/_2156_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_2900_  (.A(\wave_gen_inst/_2006_ ),
    .B(\wave_gen_inst/_2007_ ),
    .C(\wave_gen_inst/_2156_ ),
    .X(\wave_gen_inst/_2157_ ));
 sky130_fd_sc_hd__o22a_1 \wave_gen_inst/_2901_  (.A1(\wave_gen_inst/_1980_ ),
    .A2(\wave_gen_inst/_1996_ ),
    .B1(\wave_gen_inst/_2000_ ),
    .B2(\wave_gen_inst/_1995_ ),
    .X(\wave_gen_inst/_2158_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2902_  (.A(\wave_gen_inst/_2009_ ),
    .B(\wave_gen_inst/_2012_ ),
    .C(\wave_gen_inst/_2013_ ),
    .X(\wave_gen_inst/_2159_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2903_  (.A(\wave_gen_inst/param1[1] ),
    .B(net474),
    .Y(\wave_gen_inst/_2160_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_2904_  (.A(\wave_gen_inst/_1996_ ),
    .B(\wave_gen_inst/_2160_ ),
    .X(\wave_gen_inst/_2161_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2905_  (.A(\wave_gen_inst/_2159_ ),
    .B(\wave_gen_inst/_2161_ ),
    .Y(\wave_gen_inst/_2162_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2906_  (.A(\wave_gen_inst/_2158_ ),
    .B(\wave_gen_inst/_2162_ ),
    .Y(\wave_gen_inst/_2163_ ));
 sky130_fd_sc_hd__a32o_1 \wave_gen_inst/_2907_  (.A1(\wave_gen_inst/_1963_ ),
    .A2(\wave_gen_inst/_1967_ ),
    .A3(\wave_gen_inst/_2026_ ),
    .B1(\wave_gen_inst/_2027_ ),
    .B2(\wave_gen_inst/_2015_ ),
    .X(\wave_gen_inst/_2164_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2908_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_2165_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2909_  (.A(\wave_gen_inst/_2008_ ),
    .B(\wave_gen_inst/_2011_ ),
    .Y(\wave_gen_inst/_2166_ ));
 sky130_fd_sc_hd__a2bb2oi_2 \wave_gen_inst/_2910_  (.A1_N(\wave_gen_inst/_1971_ ),
    .A2_N(\wave_gen_inst/_2165_ ),
    .B1(\wave_gen_inst/_2166_ ),
    .B2(\wave_gen_inst/_2010_ ),
    .Y(\wave_gen_inst/_2167_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2911_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_2168_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2912_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_2169_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2913_  (.A(\wave_gen_inst/_2165_ ),
    .B(\wave_gen_inst/_2168_ ),
    .C(\wave_gen_inst/_2169_ ),
    .X(\wave_gen_inst/_2170_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2914_  (.A(\wave_gen_inst/_2019_ ),
    .B(\wave_gen_inst/_2020_ ),
    .C(\wave_gen_inst/_2021_ ),
    .X(\wave_gen_inst/_2171_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2915_  (.A(\wave_gen_inst/_2170_ ),
    .B(\wave_gen_inst/_2171_ ),
    .Y(\wave_gen_inst/_2172_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2916_  (.A(\wave_gen_inst/_2167_ ),
    .B(\wave_gen_inst/_2172_ ),
    .Y(\wave_gen_inst/_2173_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2917_  (.A(\wave_gen_inst/_2018_ ),
    .B(\wave_gen_inst/_2022_ ),
    .C(\wave_gen_inst/_2025_ ),
    .X(\wave_gen_inst/_2174_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2918_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_2175_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2919_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_2176_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2920_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_2177_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2921_  (.A(\wave_gen_inst/_2175_ ),
    .B(\wave_gen_inst/_2176_ ),
    .C(\wave_gen_inst/_2177_ ),
    .X(\wave_gen_inst/_2178_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_2922_  (.A(\wave_gen_inst/_2017_ ),
    .B(\wave_gen_inst/_2023_ ),
    .C(\wave_gen_inst/_2024_ ),
    .X(\wave_gen_inst/_2179_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2923_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[1] ),
    .Y(\wave_gen_inst/_2180_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2924_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_2181_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2925_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_2182_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2926_  (.A(\wave_gen_inst/_2180_ ),
    .B(\wave_gen_inst/_2181_ ),
    .C(\wave_gen_inst/_2182_ ),
    .X(\wave_gen_inst/_2183_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_2927_  (.A(\wave_gen_inst/_2178_ ),
    .B(\wave_gen_inst/_2179_ ),
    .C(\wave_gen_inst/_2183_ ),
    .X(\wave_gen_inst/_2184_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_2928_  (.A(\wave_gen_inst/_2174_ ),
    .B(\wave_gen_inst/_2184_ ),
    .X(\wave_gen_inst/_2185_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2929_  (.A(\wave_gen_inst/_2173_ ),
    .B(\wave_gen_inst/_2185_ ),
    .Y(\wave_gen_inst/_2186_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_2930_  (.A(\wave_gen_inst/_2164_ ),
    .B(\wave_gen_inst/_2186_ ),
    .X(\wave_gen_inst/_2187_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2931_  (.A(\wave_gen_inst/_2163_ ),
    .B(\wave_gen_inst/_2187_ ),
    .Y(\wave_gen_inst/_2188_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2932_  (.A(\wave_gen_inst/_2157_ ),
    .B(\wave_gen_inst/_2188_ ),
    .Y(\wave_gen_inst/_2189_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_2933_  (.A(\wave_gen_inst/_2155_ ),
    .B(\wave_gen_inst/_2189_ ),
    .Y(\wave_gen_inst/_2190_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_2934_  (.A(\wave_gen_inst/_2154_ ),
    .B(\wave_gen_inst/_2190_ ),
    .X(\wave_gen_inst/_2191_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_2935_  (.A(\wave_gen_inst/_2152_ ),
    .B(\wave_gen_inst/_2191_ ),
    .X(\wave_gen_inst/_2192_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2936_  (.A(\wave_gen_inst/_1901_ ),
    .B(\wave_gen_inst/_2192_ ),
    .Y(\wave_gen_inst/_2193_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2937_  (.A(\wave_gen_inst/_2150_ ),
    .B(\wave_gen_inst/_2058_ ),
    .C(\wave_gen_inst/_2149_ ),
    .Y(\wave_gen_inst/_2194_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \wave_gen_inst/_2938_  (.A(\wave_gen_inst/_2151_ ),
    .SLEEP(\wave_gen_inst/_2194_ ),
    .X(\wave_gen_inst/_2195_ ));
 sky130_fd_sc_hd__and3_4 \wave_gen_inst/_2946_  (.A(net13),
    .B(net11),
    .C(net12),
    .X(\wave_gen_inst/_0106_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_2948_  (.A(net163),
    .B(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_0108_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2949_  (.A1(\wave_gen_inst/_2193_ ),
    .A2(\wave_gen_inst/_2195_ ),
    .B1(\wave_gen_inst/_0108_ ),
    .Y(\wave_gen_inst/_0109_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2950_  (.A1(\wave_gen_inst/_2193_ ),
    .A2(\wave_gen_inst/_2195_ ),
    .B1(\wave_gen_inst/_0109_ ),
    .Y(\wave_gen_inst/_0110_ ));
 sky130_fd_sc_hd__nand3_4 \wave_gen_inst/_2951_  (.A(net13),
    .B(net11),
    .C(net12),
    .Y(\wave_gen_inst/_0111_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_2952_  (.A(net163),
    .B(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_0112_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2953_  (.A(\wave_gen_inst/_2192_ ),
    .B(\wave_gen_inst/_0112_ ),
    .Y(\wave_gen_inst/_0113_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2954_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/_1655_ ),
    .Y(\wave_gen_inst/_0114_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_2955_  (.A_N(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/counter[3] ),
    .Y(\wave_gen_inst/_0115_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2956_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/counter[2] ),
    .Y(\wave_gen_inst/_0116_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_2957_  (.A(\wave_gen_inst/_0114_ ),
    .B(\wave_gen_inst/_0115_ ),
    .C(\wave_gen_inst/_0116_ ),
    .Y(\wave_gen_inst/_0117_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_2958_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/counter[1] ),
    .Y(\wave_gen_inst/_0118_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_2959_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1550_ ),
    .B1(\wave_gen_inst/_0118_ ),
    .Y(\wave_gen_inst/_0119_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_2960_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/counter[1] ),
    .B1(\wave_gen_inst/_0119_ ),
    .Y(\wave_gen_inst/_0120_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_2961_  (.A_N(\wave_gen_inst/_0117_ ),
    .B(\wave_gen_inst/_0120_ ),
    .Y(\wave_gen_inst/_0121_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_2962_  (.A_N(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/_0115_ ),
    .C(\wave_gen_inst/param2[3] ),
    .Y(\wave_gen_inst/_0122_ ));
 sky130_fd_sc_hd__inv_4 \wave_gen_inst/_2963_  (.A(net846),
    .Y(\wave_gen_inst/_0123_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2964_  (.A(\wave_gen_inst/counter[11] ),
    .Y(\wave_gen_inst/_0124_ ));
 sky130_fd_sc_hd__o221a_1 \wave_gen_inst/_2965_  (.A1(\wave_gen_inst/param2[10] ),
    .A2(\wave_gen_inst/_1646_ ),
    .B1(\wave_gen_inst/_0123_ ),
    .B2(\wave_gen_inst/param2[11] ),
    .C1(\wave_gen_inst/_0124_ ),
    .X(\wave_gen_inst/_0125_ ));
 sky130_fd_sc_hd__a22oi_2 \wave_gen_inst/_2966_  (.A1(\wave_gen_inst/param2[9] ),
    .A2(\wave_gen_inst/_1590_ ),
    .B1(\wave_gen_inst/_1646_ ),
    .B2(\wave_gen_inst/param2[10] ),
    .Y(\wave_gen_inst/_0126_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2967_  (.A(\wave_gen_inst/param2[11] ),
    .B(\wave_gen_inst/_0123_ ),
    .Y(\wave_gen_inst/_0127_ ));
 sky130_fd_sc_hd__o2111ai_2 \wave_gen_inst/_2968_  (.A1(\wave_gen_inst/param2[9] ),
    .A2(\wave_gen_inst/_1590_ ),
    .B1(\wave_gen_inst/_0125_ ),
    .C1(\wave_gen_inst/_0126_ ),
    .D1(\wave_gen_inst/_0127_ ),
    .Y(\wave_gen_inst/_0128_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_2969_  (.A(\wave_gen_inst/param2[5] ),
    .SLEEP(\wave_gen_inst/counter[4] ),
    .X(\wave_gen_inst/_0129_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_2970_  (.A(\wave_gen_inst/param2[6] ),
    .Y(\wave_gen_inst/_0130_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_2971_  (.A1(\wave_gen_inst/param2[5] ),
    .A2(\wave_gen_inst/_1578_ ),
    .B1(\wave_gen_inst/counter[5] ),
    .B2(\wave_gen_inst/_0130_ ),
    .Y(\wave_gen_inst/_0131_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2972_  (.A1(\wave_gen_inst/_0130_ ),
    .A2(\wave_gen_inst/counter[5] ),
    .B1(\wave_gen_inst/_0131_ ),
    .Y(\wave_gen_inst/_0132_ ));
 sky130_fd_sc_hd__clkinv_4 \wave_gen_inst/_2973_  (.A(\wave_gen_inst/counter[7] ),
    .Y(\wave_gen_inst/_0133_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_2974_  (.A(\wave_gen_inst/param2[7] ),
    .SLEEP(\wave_gen_inst/counter[6] ),
    .X(\wave_gen_inst/_0134_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2975_  (.A(\wave_gen_inst/counter[6] ),
    .Y(\wave_gen_inst/_0135_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_2976_  (.A1(\wave_gen_inst/param2[7] ),
    .A2(\wave_gen_inst/_0135_ ),
    .B1(\wave_gen_inst/_0133_ ),
    .B2(\wave_gen_inst/param2[8] ),
    .Y(\wave_gen_inst/_0136_ ));
 sky130_fd_sc_hd__a211oi_2 \wave_gen_inst/_2977_  (.A1(\wave_gen_inst/param2[8] ),
    .A2(\wave_gen_inst/_0133_ ),
    .B1(\wave_gen_inst/_0134_ ),
    .C1(\wave_gen_inst/_0136_ ),
    .Y(\wave_gen_inst/_0137_ ));
 sky130_fd_sc_hd__nand4bb_2 \wave_gen_inst/_2978_  (.A_N(\wave_gen_inst/_0128_ ),
    .B_N(\wave_gen_inst/_0129_ ),
    .C(\wave_gen_inst/_0132_ ),
    .D(\wave_gen_inst/_0137_ ),
    .Y(\wave_gen_inst/_0138_ ));
 sky130_fd_sc_hd__a31oi_2 \wave_gen_inst/_2979_  (.A1(\wave_gen_inst/_0114_ ),
    .A2(\wave_gen_inst/_0121_ ),
    .A3(\wave_gen_inst/_0122_ ),
    .B1(\wave_gen_inst/_0138_ ),
    .Y(\wave_gen_inst/_0139_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_2980_  (.A(\wave_gen_inst/_0125_ ),
    .SLEEP(\wave_gen_inst/_0126_ ),
    .X(\wave_gen_inst/_0140_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/_2981_  (.A(\wave_gen_inst/counter[5] ),
    .Y(\wave_gen_inst/_0141_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2982_  (.A1(\wave_gen_inst/param2[6] ),
    .A2(\wave_gen_inst/_0141_ ),
    .B1(\wave_gen_inst/_0129_ ),
    .Y(\wave_gen_inst/_0142_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2983_  (.A1(\wave_gen_inst/_0130_ ),
    .A2(\wave_gen_inst/counter[5] ),
    .B1(\wave_gen_inst/_0142_ ),
    .Y(\wave_gen_inst/_0143_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_2984_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/_0133_ ),
    .C(\wave_gen_inst/_0134_ ),
    .X(\wave_gen_inst/_0144_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_2985_  (.A1(\wave_gen_inst/_0137_ ),
    .A2(\wave_gen_inst/_0143_ ),
    .B1(\wave_gen_inst/_0144_ ),
    .Y(\wave_gen_inst/_0145_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_2986_  (.A1(\wave_gen_inst/counter[11] ),
    .A2(\wave_gen_inst/_0127_ ),
    .B1(\wave_gen_inst/_0128_ ),
    .B2(\wave_gen_inst/_0145_ ),
    .Y(\wave_gen_inst/_0146_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2987_  (.A(\wave_gen_inst/_0139_ ),
    .B(\wave_gen_inst/_0140_ ),
    .C(\wave_gen_inst/_0146_ ),
    .Y(\wave_gen_inst/_0147_ ));
 sky130_fd_sc_hd__a2111oi_4 \wave_gen_inst/_2988_  (.A1(\wave_gen_inst/param2[1] ),
    .A2(\wave_gen_inst/_1550_ ),
    .B1(\wave_gen_inst/_0138_ ),
    .C1(\wave_gen_inst/_0117_ ),
    .D1(\wave_gen_inst/_0119_ ),
    .Y(\wave_gen_inst/_0148_ ));
 sky130_fd_sc_hd__or3_2 \wave_gen_inst/_2989_  (.A(\wave_gen_inst/counter[13] ),
    .B(\wave_gen_inst/counter[14] ),
    .C(\wave_gen_inst/counter[15] ),
    .X(\wave_gen_inst/_0149_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2991_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/counter[25] ),
    .Y(\wave_gen_inst/_0151_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_2992_  (.A(\wave_gen_inst/counter[30] ),
    .B(\wave_gen_inst/counter[31] ),
    .Y(\wave_gen_inst/_0152_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2993_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/counter[21] ),
    .C(\wave_gen_inst/counter[22] ),
    .Y(\wave_gen_inst/_0153_ ));
 sky130_fd_sc_hd__or2_2 \wave_gen_inst/_2994_  (.A(\wave_gen_inst/counter[17] ),
    .B(\wave_gen_inst/counter[18] ),
    .X(\wave_gen_inst/_0154_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_2995_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/counter[19] ),
    .C(\wave_gen_inst/_0154_ ),
    .Y(\wave_gen_inst/_0155_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_2996_  (.A(\wave_gen_inst/_0153_ ),
    .B(\wave_gen_inst/_0155_ ),
    .Y(\wave_gen_inst/_0156_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_2997_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_0156_ ),
    .Y(\wave_gen_inst/_0157_ ));
 sky130_fd_sc_hd__nor4_2 \wave_gen_inst/_2999_  (.A(\wave_gen_inst/counter[26] ),
    .B(\wave_gen_inst/counter[27] ),
    .C(\wave_gen_inst/counter[28] ),
    .D(\wave_gen_inst/counter[29] ),
    .Y(\wave_gen_inst/_0159_ ));
 sky130_fd_sc_hd__nand4_4 \wave_gen_inst/_3000_  (.A(\wave_gen_inst/_0151_ ),
    .B(\wave_gen_inst/_0152_ ),
    .C(\wave_gen_inst/_0157_ ),
    .D(\wave_gen_inst/_0159_ ),
    .Y(\wave_gen_inst/_0160_ ));
 sky130_fd_sc_hd__nor3_4 \wave_gen_inst/_3001_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/_0149_ ),
    .C(\wave_gen_inst/_0160_ ),
    .Y(\wave_gen_inst/_0161_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_3002_  (.A(net11),
    .B(net12),
    .Y(\wave_gen_inst/_0162_ ));
 sky130_fd_sc_hd__nand3_2 \wave_gen_inst/_3003_  (.A(net13),
    .B(\wave_gen_inst/_0161_ ),
    .C(\wave_gen_inst/_0162_ ),
    .Y(\wave_gen_inst/_0163_ ));
 sky130_fd_sc_hd__nor3_4 \wave_gen_inst/_3004_  (.A(\wave_gen_inst/_0147_ ),
    .B(\wave_gen_inst/_0148_ ),
    .C(\wave_gen_inst/_0163_ ),
    .Y(\wave_gen_inst/_0164_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_3006_  (.A1(net11),
    .A2(net12),
    .B1(net13),
    .Y(\wave_gen_inst/_0166_ ));
 sky130_fd_sc_hd__a21oi_4 \wave_gen_inst/_3007_  (.A1(net11),
    .A2(net12),
    .B1(\wave_gen_inst/_0166_ ),
    .Y(\wave_gen_inst/_0167_ ));
 sky130_fd_sc_hd__nor2_8 \wave_gen_inst/_3009_  (.A(net13),
    .B(\wave_gen_inst/_0162_ ),
    .Y(\wave_gen_inst/_0169_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3011_  (.A1(\wave_gen_inst/param1[1] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[1] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net26),
    .Y(\wave_gen_inst/_0171_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3013_  (.A1(\wave_gen_inst/_0110_ ),
    .A2(\wave_gen_inst/_0113_ ),
    .A3(\wave_gen_inst/_0171_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0000_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3015_  (.A(\wave_gen_inst/_1901_ ),
    .B(\wave_gen_inst/_2192_ ),
    .C(\wave_gen_inst/_2195_ ),
    .X(\wave_gen_inst/_0174_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3016_  (.A(\wave_gen_inst/_2154_ ),
    .B(\wave_gen_inst/_2190_ ),
    .Y(\wave_gen_inst/_0175_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/_3017_  (.A1(\wave_gen_inst/_2033_ ),
    .A2(\wave_gen_inst/_2151_ ),
    .B1_N(\wave_gen_inst/_2191_ ),
    .Y(\wave_gen_inst/_0176_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3018_  (.A(\wave_gen_inst/_2155_ ),
    .B(\wave_gen_inst/_2189_ ),
    .Y(\wave_gen_inst/_0177_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3019_  (.A1(\wave_gen_inst/_2157_ ),
    .A2(\wave_gen_inst/_2188_ ),
    .B1(\wave_gen_inst/_0177_ ),
    .Y(\wave_gen_inst/_0178_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3020_  (.A(\wave_gen_inst/_2161_ ),
    .Y(\wave_gen_inst/_0179_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3021_  (.A(\wave_gen_inst/_2158_ ),
    .B(\wave_gen_inst/_2159_ ),
    .C(\wave_gen_inst/_0179_ ),
    .X(\wave_gen_inst/_0180_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3022_  (.A(\wave_gen_inst/_2164_ ),
    .SLEEP(\wave_gen_inst/_2186_ ),
    .X(\wave_gen_inst/_0181_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3023_  (.A(\wave_gen_inst/_2163_ ),
    .SLEEP(\wave_gen_inst/_2187_ ),
    .X(\wave_gen_inst/_0182_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3024_  (.A(\wave_gen_inst/_0181_ ),
    .B(\wave_gen_inst/_0182_ ),
    .Y(\wave_gen_inst/_0183_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3025_  (.A(\wave_gen_inst/_2174_ ),
    .B(\wave_gen_inst/_2184_ ),
    .X(\wave_gen_inst/_0184_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3026_  (.A1(\wave_gen_inst/_2173_ ),
    .A2(\wave_gen_inst/_2185_ ),
    .B1(\wave_gen_inst/_0184_ ),
    .Y(\wave_gen_inst/_0185_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3027_  (.A(\wave_gen_inst/_2165_ ),
    .B(\wave_gen_inst/_2168_ ),
    .C(\wave_gen_inst/_2169_ ),
    .X(\wave_gen_inst/_0186_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3028_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0187_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3029_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0188_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3030_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0189_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3031_  (.A(\wave_gen_inst/_0188_ ),
    .B(\wave_gen_inst/_0189_ ),
    .X(\wave_gen_inst/_0190_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3032_  (.A(\wave_gen_inst/_0187_ ),
    .B(\wave_gen_inst/_0190_ ),
    .Y(\wave_gen_inst/_0191_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3033_  (.A(\wave_gen_inst/_2175_ ),
    .B(\wave_gen_inst/_2176_ ),
    .C(\wave_gen_inst/_2177_ ),
    .X(\wave_gen_inst/_0192_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3034_  (.A(\wave_gen_inst/_0191_ ),
    .B(\wave_gen_inst/_0192_ ),
    .X(\wave_gen_inst/_0193_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3035_  (.A(\wave_gen_inst/_0186_ ),
    .B(\wave_gen_inst/_0193_ ),
    .X(\wave_gen_inst/_0194_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3036_  (.A(\wave_gen_inst/_2179_ ),
    .B(\wave_gen_inst/_2183_ ),
    .Y(\wave_gen_inst/_0195_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3037_  (.A_N(\wave_gen_inst/_2179_ ),
    .B(\wave_gen_inst/_2183_ ),
    .Y(\wave_gen_inst/_0196_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/_3038_  (.A1(\wave_gen_inst/_2178_ ),
    .A2(\wave_gen_inst/_0195_ ),
    .B1_N(\wave_gen_inst/_0196_ ),
    .Y(\wave_gen_inst/_0197_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3039_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_0198_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3040_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_0199_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3041_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_0200_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3042_  (.A(\wave_gen_inst/_0199_ ),
    .B(\wave_gen_inst/_0200_ ),
    .X(\wave_gen_inst/_0201_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3043_  (.A(\wave_gen_inst/_0198_ ),
    .B(\wave_gen_inst/_0201_ ),
    .Y(\wave_gen_inst/_0202_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3044_  (.A(\wave_gen_inst/_2180_ ),
    .B(\wave_gen_inst/_2181_ ),
    .C(\wave_gen_inst/_2182_ ),
    .X(\wave_gen_inst/_0203_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3045_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[2] ),
    .Y(\wave_gen_inst/_0204_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3046_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_0205_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3047_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_0206_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_3048_  (.A(\wave_gen_inst/_0204_ ),
    .B(\wave_gen_inst/_0205_ ),
    .C(\wave_gen_inst/_0206_ ),
    .X(\wave_gen_inst/_0207_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3049_  (.A(\wave_gen_inst/_0203_ ),
    .B(\wave_gen_inst/_0207_ ),
    .Y(\wave_gen_inst/_0208_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3050_  (.A(\wave_gen_inst/_0202_ ),
    .B(\wave_gen_inst/_0208_ ),
    .X(\wave_gen_inst/_0209_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3051_  (.A(\wave_gen_inst/_0197_ ),
    .B(\wave_gen_inst/_0209_ ),
    .Y(\wave_gen_inst/_0210_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3052_  (.A(\wave_gen_inst/_0194_ ),
    .B(\wave_gen_inst/_0210_ ),
    .Y(\wave_gen_inst/_0211_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3053_  (.A(\wave_gen_inst/_0185_ ),
    .B(\wave_gen_inst/_0211_ ),
    .X(\wave_gen_inst/_0212_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3054_  (.A(\wave_gen_inst/_2170_ ),
    .Y(\wave_gen_inst/_0213_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_3055_  (.A(\wave_gen_inst/_2167_ ),
    .B(\wave_gen_inst/_0213_ ),
    .C(\wave_gen_inst/_2171_ ),
    .X(\wave_gen_inst/_0214_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3056_  (.A(\wave_gen_inst/param1[2] ),
    .B(net475),
    .C(\wave_gen_inst/_1998_ ),
    .Y(\wave_gen_inst/_0215_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3057_  (.A(\wave_gen_inst/_0214_ ),
    .B(\wave_gen_inst/_0215_ ),
    .X(\wave_gen_inst/_0216_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3058_  (.A(\wave_gen_inst/_0212_ ),
    .B(\wave_gen_inst/_0216_ ),
    .X(\wave_gen_inst/_0217_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3059_  (.A(\wave_gen_inst/_0183_ ),
    .B(\wave_gen_inst/_0217_ ),
    .X(\wave_gen_inst/_0218_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3060_  (.A(\wave_gen_inst/_0180_ ),
    .B(\wave_gen_inst/_0218_ ),
    .Y(\wave_gen_inst/_0219_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3061_  (.A(\wave_gen_inst/_0178_ ),
    .B(\wave_gen_inst/_0219_ ),
    .X(\wave_gen_inst/_0220_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3062_  (.A1(\wave_gen_inst/_0175_ ),
    .A2(\wave_gen_inst/_0176_ ),
    .B1(\wave_gen_inst/_0220_ ),
    .X(\wave_gen_inst/_0221_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3063_  (.A(\wave_gen_inst/_0175_ ),
    .B(\wave_gen_inst/_0176_ ),
    .C(\wave_gen_inst/_0220_ ),
    .Y(\wave_gen_inst/_0222_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3064_  (.A(\wave_gen_inst/_0221_ ),
    .B(\wave_gen_inst/_0222_ ),
    .Y(\wave_gen_inst/_0223_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3065_  (.A(\wave_gen_inst/_1814_ ),
    .B(\wave_gen_inst/_0223_ ),
    .Y(\wave_gen_inst/_0224_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3066_  (.A(\wave_gen_inst/_0174_ ),
    .B(\wave_gen_inst/_0224_ ),
    .Y(\wave_gen_inst/_0225_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3067_  (.A(\wave_gen_inst/_0174_ ),
    .B(\wave_gen_inst/_0224_ ),
    .Y(\wave_gen_inst/_0226_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3068_  (.A(\wave_gen_inst/_0108_ ),
    .B(\wave_gen_inst/_0226_ ),
    .Y(\wave_gen_inst/_0227_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3069_  (.A(\wave_gen_inst/_0112_ ),
    .B(\wave_gen_inst/_0223_ ),
    .Y(\wave_gen_inst/_0228_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3070_  (.A1(\wave_gen_inst/param1[2] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[2] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net37),
    .Y(\wave_gen_inst/_0229_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3071_  (.A(\wave_gen_inst/_0228_ ),
    .B(\wave_gen_inst/_0229_ ),
    .Y(\wave_gen_inst/_0230_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3072_  (.A1(\wave_gen_inst/_0225_ ),
    .A2(\wave_gen_inst/_0227_ ),
    .B1(\wave_gen_inst/_0230_ ),
    .Y(\wave_gen_inst/_0231_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3073_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0231_ ),
    .Y(\wave_gen_inst/_0001_ ));
 sky130_fd_sc_hd__inv_8 \wave_gen_inst/_3074_  (.A(net162),
    .Y(\wave_gen_inst/_0232_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_3075_  (.A(\wave_gen_inst/_0232_ ),
    .B(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_0233_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3076_  (.A(\wave_gen_inst/_1814_ ),
    .B(\wave_gen_inst/_0174_ ),
    .C(\wave_gen_inst/_0223_ ),
    .X(\wave_gen_inst/_0234_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3077_  (.A(\wave_gen_inst/_0178_ ),
    .B(\wave_gen_inst/_0219_ ),
    .Y(\wave_gen_inst/_0235_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3078_  (.A(\wave_gen_inst/_0217_ ),
    .SLEEP(\wave_gen_inst/_0183_ ),
    .X(\wave_gen_inst/_0236_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3079_  (.A(\wave_gen_inst/_0180_ ),
    .B(\wave_gen_inst/_0218_ ),
    .Y(\wave_gen_inst/_0237_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3080_  (.A(\wave_gen_inst/_0236_ ),
    .B(\wave_gen_inst/_0237_ ),
    .Y(\wave_gen_inst/_0238_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3081_  (.A(\wave_gen_inst/_0185_ ),
    .B(\wave_gen_inst/_0211_ ),
    .Y(\wave_gen_inst/_0239_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3082_  (.A1(\wave_gen_inst/_0212_ ),
    .A2(\wave_gen_inst/_0216_ ),
    .B1(\wave_gen_inst/_0239_ ),
    .Y(\wave_gen_inst/_0240_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3083_  (.A(\wave_gen_inst/_0191_ ),
    .SLEEP(\wave_gen_inst/_0192_ ),
    .X(\wave_gen_inst/_0241_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3084_  (.A(\wave_gen_inst/_0186_ ),
    .B(\wave_gen_inst/_0193_ ),
    .Y(\wave_gen_inst/_0242_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3085_  (.A(\wave_gen_inst/_0241_ ),
    .B(\wave_gen_inst/_0242_ ),
    .Y(\wave_gen_inst/_0243_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3086_  (.A(\wave_gen_inst/_0209_ ),
    .SLEEP(\wave_gen_inst/_0197_ ),
    .X(\wave_gen_inst/_0244_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3087_  (.A1(\wave_gen_inst/_0194_ ),
    .A2(\wave_gen_inst/_0210_ ),
    .B1(\wave_gen_inst/_0244_ ),
    .Y(\wave_gen_inst/_0245_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3088_  (.A(\wave_gen_inst/_0188_ ),
    .B(\wave_gen_inst/_0187_ ),
    .C(\wave_gen_inst/_0189_ ),
    .X(\wave_gen_inst/_0246_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3089_  (.A(\wave_gen_inst/param1[3] ),
    .B(net476),
    .Y(\wave_gen_inst/_0247_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3090_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0248_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3092_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0250_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3093_  (.A(\wave_gen_inst/_0248_ ),
    .B(\wave_gen_inst/_0250_ ),
    .X(\wave_gen_inst/_0251_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3094_  (.A(\wave_gen_inst/_0247_ ),
    .B(\wave_gen_inst/_0251_ ),
    .Y(\wave_gen_inst/_0252_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3095_  (.A(\wave_gen_inst/_0199_ ),
    .B(\wave_gen_inst/_0198_ ),
    .C(\wave_gen_inst/_0200_ ),
    .X(\wave_gen_inst/_0253_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3096_  (.A(\wave_gen_inst/_0252_ ),
    .B(\wave_gen_inst/_0253_ ),
    .X(\wave_gen_inst/_0254_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3097_  (.A(\wave_gen_inst/_0246_ ),
    .B(\wave_gen_inst/_0254_ ),
    .X(\wave_gen_inst/_0255_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3098_  (.A(\wave_gen_inst/_0207_ ),
    .SLEEP(\wave_gen_inst/_0203_ ),
    .X(\wave_gen_inst/_0256_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3099_  (.A1(\wave_gen_inst/_0202_ ),
    .A2(\wave_gen_inst/_0208_ ),
    .B1(\wave_gen_inst/_0256_ ),
    .Y(\wave_gen_inst/_0257_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3100_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0258_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3101_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_0259_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3102_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_0260_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3103_  (.A(\wave_gen_inst/_0259_ ),
    .B(\wave_gen_inst/_0260_ ),
    .X(\wave_gen_inst/_0261_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3104_  (.A(\wave_gen_inst/_0258_ ),
    .B(\wave_gen_inst/_0261_ ),
    .Y(\wave_gen_inst/_0262_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3105_  (.A(\wave_gen_inst/_0204_ ),
    .B(\wave_gen_inst/_0205_ ),
    .C(\wave_gen_inst/_0206_ ),
    .X(\wave_gen_inst/_0263_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3106_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_0264_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3107_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[3] ),
    .Y(\wave_gen_inst/_0265_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3108_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_0266_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3109_  (.A(\wave_gen_inst/_0265_ ),
    .B(\wave_gen_inst/_0266_ ),
    .X(\wave_gen_inst/_0267_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3110_  (.A(\wave_gen_inst/_0264_ ),
    .B(\wave_gen_inst/_0267_ ),
    .Y(\wave_gen_inst/_0268_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3111_  (.A(\wave_gen_inst/_0263_ ),
    .B(\wave_gen_inst/_0268_ ),
    .Y(\wave_gen_inst/_0269_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3112_  (.A(\wave_gen_inst/_0262_ ),
    .B(\wave_gen_inst/_0269_ ),
    .X(\wave_gen_inst/_0270_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3113_  (.A(\wave_gen_inst/_0257_ ),
    .B(\wave_gen_inst/_0270_ ),
    .Y(\wave_gen_inst/_0271_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3114_  (.A(\wave_gen_inst/_0255_ ),
    .B(\wave_gen_inst/_0271_ ),
    .Y(\wave_gen_inst/_0272_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3115_  (.A(\wave_gen_inst/_0245_ ),
    .B(\wave_gen_inst/_0272_ ),
    .Y(\wave_gen_inst/_0273_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3116_  (.A(\wave_gen_inst/_0243_ ),
    .B(\wave_gen_inst/_0273_ ),
    .Y(\wave_gen_inst/_0274_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3117_  (.A(\wave_gen_inst/_0240_ ),
    .B(\wave_gen_inst/_0274_ ),
    .X(\wave_gen_inst/_0275_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3119_  (.A(\wave_gen_inst/_1998_ ),
    .B(\wave_gen_inst/_0214_ ),
    .Y(\wave_gen_inst/_0277_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3120_  (.A(\wave_gen_inst/param1[2] ),
    .B(net477),
    .C(\wave_gen_inst/_0277_ ),
    .Y(\wave_gen_inst/_0278_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3121_  (.A(\wave_gen_inst/_0275_ ),
    .B(\wave_gen_inst/_0278_ ),
    .Y(\wave_gen_inst/_0279_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3122_  (.A(\wave_gen_inst/_0238_ ),
    .B(\wave_gen_inst/_0279_ ),
    .Y(\wave_gen_inst/_0280_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3123_  (.A1(\wave_gen_inst/_0235_ ),
    .A2(\wave_gen_inst/_0221_ ),
    .B1(\wave_gen_inst/_0280_ ),
    .X(\wave_gen_inst/_0281_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3124_  (.A(\wave_gen_inst/_0235_ ),
    .B(\wave_gen_inst/_0221_ ),
    .C(\wave_gen_inst/_0280_ ),
    .Y(\wave_gen_inst/_0282_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3125_  (.A(\wave_gen_inst/_0281_ ),
    .B(\wave_gen_inst/_0282_ ),
    .Y(\wave_gen_inst/_0283_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3126_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/_0283_ ),
    .Y(\wave_gen_inst/_0284_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3127_  (.A(\wave_gen_inst/_0234_ ),
    .B(\wave_gen_inst/_0284_ ),
    .Y(\wave_gen_inst/_0285_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3128_  (.A(\wave_gen_inst/_0233_ ),
    .B(\wave_gen_inst/_0285_ ),
    .Y(\wave_gen_inst/_0286_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3129_  (.A(\wave_gen_inst/_0112_ ),
    .B(\wave_gen_inst/_0283_ ),
    .Y(\wave_gen_inst/_0287_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3130_  (.A1(\wave_gen_inst/param1[3] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[3] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net40),
    .Y(\wave_gen_inst/_0288_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3131_  (.A1(\wave_gen_inst/_0286_ ),
    .A2(\wave_gen_inst/_0287_ ),
    .A3(\wave_gen_inst/_0288_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0002_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3132_  (.A1(\wave_gen_inst/_0236_ ),
    .A2(\wave_gen_inst/_0237_ ),
    .B1(\wave_gen_inst/_0279_ ),
    .Y(\wave_gen_inst/_0289_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3133_  (.A(\wave_gen_inst/_0289_ ),
    .Y(\wave_gen_inst/_0290_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3134_  (.A(\wave_gen_inst/_0290_ ),
    .B(\wave_gen_inst/_0281_ ),
    .Y(\wave_gen_inst/_0291_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3135_  (.A(\wave_gen_inst/_0240_ ),
    .B(\wave_gen_inst/_0274_ ),
    .C(\wave_gen_inst/_0278_ ),
    .X(\wave_gen_inst/_0292_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3136_  (.A(\wave_gen_inst/_0243_ ),
    .B(\wave_gen_inst/_0245_ ),
    .C(\wave_gen_inst/_0272_ ),
    .X(\wave_gen_inst/_0293_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3137_  (.A(\wave_gen_inst/_0252_ ),
    .SLEEP(\wave_gen_inst/_0253_ ),
    .X(\wave_gen_inst/_0294_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3138_  (.A(\wave_gen_inst/_0246_ ),
    .B(\wave_gen_inst/_0254_ ),
    .Y(\wave_gen_inst/_0295_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3139_  (.A(\wave_gen_inst/_0294_ ),
    .B(\wave_gen_inst/_0295_ ),
    .Y(\wave_gen_inst/_0296_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3140_  (.A_N(\wave_gen_inst/_0257_ ),
    .B(\wave_gen_inst/_0270_ ),
    .Y(\wave_gen_inst/_0297_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/_3141_  (.A1(\wave_gen_inst/_0255_ ),
    .A2(\wave_gen_inst/_0271_ ),
    .B1_N(\wave_gen_inst/_0297_ ),
    .Y(\wave_gen_inst/_0298_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3142_  (.A(\wave_gen_inst/_0248_ ),
    .B(\wave_gen_inst/_0247_ ),
    .C(\wave_gen_inst/_0250_ ),
    .X(\wave_gen_inst/_0299_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3143_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0300_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3144_  (.A(\wave_gen_inst/param1[4] ),
    .B(net478),
    .Y(\wave_gen_inst/_0301_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3145_  (.A(\wave_gen_inst/_0300_ ),
    .B(\wave_gen_inst/_0301_ ),
    .X(\wave_gen_inst/_0302_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3146_  (.A(\wave_gen_inst/_0259_ ),
    .B(\wave_gen_inst/_0258_ ),
    .C(\wave_gen_inst/_0260_ ),
    .X(\wave_gen_inst/_0303_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3147_  (.A(\wave_gen_inst/_0302_ ),
    .B(\wave_gen_inst/_0303_ ),
    .Y(\wave_gen_inst/_0304_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3148_  (.A(\wave_gen_inst/_0299_ ),
    .B(\wave_gen_inst/_0304_ ),
    .Y(\wave_gen_inst/_0305_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3149_  (.A(\wave_gen_inst/_0268_ ),
    .SLEEP(\wave_gen_inst/_0263_ ),
    .X(\wave_gen_inst/_0306_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3150_  (.A1(\wave_gen_inst/_0262_ ),
    .A2(\wave_gen_inst/_0269_ ),
    .B1(\wave_gen_inst/_0306_ ),
    .Y(\wave_gen_inst/_0307_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3151_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0308_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3152_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_0309_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3153_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0310_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3154_  (.A(\wave_gen_inst/_0309_ ),
    .B(\wave_gen_inst/_0310_ ),
    .X(\wave_gen_inst/_0311_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3155_  (.A(\wave_gen_inst/_0308_ ),
    .B(\wave_gen_inst/_0311_ ),
    .Y(\wave_gen_inst/_0312_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3156_  (.A(\wave_gen_inst/_0265_ ),
    .B(\wave_gen_inst/_0264_ ),
    .C(\wave_gen_inst/_0266_ ),
    .X(\wave_gen_inst/_0313_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3157_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_0314_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3158_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[4] ),
    .Y(\wave_gen_inst/_0315_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3159_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_0316_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3160_  (.A(\wave_gen_inst/_0315_ ),
    .B(\wave_gen_inst/_0316_ ),
    .X(\wave_gen_inst/_0317_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3161_  (.A(\wave_gen_inst/_0314_ ),
    .B(\wave_gen_inst/_0317_ ),
    .Y(\wave_gen_inst/_0318_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3162_  (.A(\wave_gen_inst/_0313_ ),
    .B(\wave_gen_inst/_0318_ ),
    .Y(\wave_gen_inst/_0319_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3163_  (.A(\wave_gen_inst/_0312_ ),
    .B(\wave_gen_inst/_0319_ ),
    .X(\wave_gen_inst/_0320_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3164_  (.A(\wave_gen_inst/_0307_ ),
    .B(\wave_gen_inst/_0320_ ),
    .Y(\wave_gen_inst/_0321_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3165_  (.A(\wave_gen_inst/_0305_ ),
    .B(\wave_gen_inst/_0321_ ),
    .Y(\wave_gen_inst/_0322_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/_3166_  (.A(\wave_gen_inst/_0296_ ),
    .B(\wave_gen_inst/_0298_ ),
    .C(\wave_gen_inst/_0322_ ),
    .X(\wave_gen_inst/_0323_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3167_  (.A(\wave_gen_inst/_0293_ ),
    .B(\wave_gen_inst/_0323_ ),
    .Y(\wave_gen_inst/_0324_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3168_  (.A(\wave_gen_inst/_0292_ ),
    .B(\wave_gen_inst/_0324_ ),
    .X(\wave_gen_inst/_0325_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_3169_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/_0291_ ),
    .C(\wave_gen_inst/_0325_ ),
    .X(\wave_gen_inst/_0326_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3170_  (.A(\wave_gen_inst/_1816_ ),
    .B(\wave_gen_inst/_0234_ ),
    .C(\wave_gen_inst/_0283_ ),
    .X(\wave_gen_inst/_0327_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3171_  (.A1(\wave_gen_inst/_0326_ ),
    .A2(\wave_gen_inst/_0327_ ),
    .B1(\wave_gen_inst/_0108_ ),
    .Y(\wave_gen_inst/_0328_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3172_  (.A1(\wave_gen_inst/_0326_ ),
    .A2(\wave_gen_inst/_0327_ ),
    .B1(\wave_gen_inst/_0328_ ),
    .Y(\wave_gen_inst/_0329_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3173_  (.A(\wave_gen_inst/_0290_ ),
    .B(\wave_gen_inst/_0281_ ),
    .C(\wave_gen_inst/_0325_ ),
    .Y(\wave_gen_inst/_0330_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_3174_  (.A1(\wave_gen_inst/_0290_ ),
    .A2(\wave_gen_inst/_0281_ ),
    .B1(\wave_gen_inst/_0325_ ),
    .Y(\wave_gen_inst/_0331_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_3175_  (.A_N(\wave_gen_inst/_0330_ ),
    .B(\wave_gen_inst/_0112_ ),
    .C(\wave_gen_inst/_0331_ ),
    .Y(\wave_gen_inst/_0332_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3176_  (.A1(\wave_gen_inst/param1[4] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[4] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net41),
    .Y(\wave_gen_inst/_0333_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3177_  (.A1(\wave_gen_inst/_0329_ ),
    .A2(\wave_gen_inst/_0332_ ),
    .A3(\wave_gen_inst/_0333_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0003_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3178_  (.A1(\wave_gen_inst/_0290_ ),
    .A2(\wave_gen_inst/_0281_ ),
    .B1(\wave_gen_inst/_0325_ ),
    .X(\wave_gen_inst/_0334_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3179_  (.A1(\wave_gen_inst/_0334_ ),
    .A2(\wave_gen_inst/_0330_ ),
    .B1(\wave_gen_inst/param1[3] ),
    .Y(\wave_gen_inst/_0335_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_3180_  (.A1(\wave_gen_inst/_0326_ ),
    .A2(\wave_gen_inst/_0327_ ),
    .B1(\wave_gen_inst/_0335_ ),
    .Y(\wave_gen_inst/_0336_ ));
 sky130_fd_sc_hd__or2_0 \wave_gen_inst/_3181_  (.A(\wave_gen_inst/_0292_ ),
    .B(\wave_gen_inst/_0324_ ),
    .X(\wave_gen_inst/_0337_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3182_  (.A(\wave_gen_inst/_0293_ ),
    .B(\wave_gen_inst/_0323_ ),
    .Y(\wave_gen_inst/_0338_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3183_  (.A(\wave_gen_inst/_0296_ ),
    .B(\wave_gen_inst/_0298_ ),
    .C(\wave_gen_inst/_0322_ ),
    .X(\wave_gen_inst/_0339_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3184_  (.A(\wave_gen_inst/_0302_ ),
    .Y(\wave_gen_inst/_0340_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3185_  (.A(\wave_gen_inst/_0299_ ),
    .B(\wave_gen_inst/_0340_ ),
    .C(\wave_gen_inst/_0303_ ),
    .X(\wave_gen_inst/_0341_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3186_  (.A_N(\wave_gen_inst/_0307_ ),
    .B(\wave_gen_inst/_0320_ ),
    .Y(\wave_gen_inst/_0342_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/_3187_  (.A1(\wave_gen_inst/_0305_ ),
    .A2(\wave_gen_inst/_0321_ ),
    .B1_N(\wave_gen_inst/_0342_ ),
    .Y(\wave_gen_inst/_0343_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3188_  (.A(\wave_gen_inst/_0318_ ),
    .SLEEP(\wave_gen_inst/_0313_ ),
    .X(\wave_gen_inst/_0344_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_3189_  (.A1(\wave_gen_inst/_0312_ ),
    .A2(\wave_gen_inst/_0319_ ),
    .B1(\wave_gen_inst/_0344_ ),
    .X(\wave_gen_inst/_0345_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3190_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0346_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3191_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0347_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3192_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0348_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3193_  (.A(\wave_gen_inst/_0347_ ),
    .B(\wave_gen_inst/_0348_ ),
    .X(\wave_gen_inst/_0349_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3194_  (.A(\wave_gen_inst/_0346_ ),
    .B(\wave_gen_inst/_0349_ ),
    .Y(\wave_gen_inst/_0350_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3195_  (.A(\wave_gen_inst/_0315_ ),
    .B(\wave_gen_inst/_0314_ ),
    .C(\wave_gen_inst/_0316_ ),
    .X(\wave_gen_inst/_0351_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3196_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_0352_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3197_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[5] ),
    .Y(\wave_gen_inst/_0353_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3198_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_0354_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3199_  (.A(\wave_gen_inst/_0353_ ),
    .B(\wave_gen_inst/_0354_ ),
    .X(\wave_gen_inst/_0355_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3200_  (.A(\wave_gen_inst/_0352_ ),
    .B(\wave_gen_inst/_0355_ ),
    .Y(\wave_gen_inst/_0356_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3201_  (.A(\wave_gen_inst/_0351_ ),
    .B(\wave_gen_inst/_0356_ ),
    .Y(\wave_gen_inst/_0357_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3202_  (.A(\wave_gen_inst/_0350_ ),
    .B(\wave_gen_inst/_0357_ ),
    .X(\wave_gen_inst/_0358_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3203_  (.A(\wave_gen_inst/_0345_ ),
    .B(\wave_gen_inst/_0358_ ),
    .Y(\wave_gen_inst/_0359_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3204_  (.A(\wave_gen_inst/_0309_ ),
    .B(\wave_gen_inst/_0308_ ),
    .C(\wave_gen_inst/_0310_ ),
    .X(\wave_gen_inst/_0360_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3205_  (.A(\wave_gen_inst/param1[5] ),
    .B(net479),
    .C(\wave_gen_inst/_0250_ ),
    .Y(\wave_gen_inst/_0361_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3206_  (.A(\wave_gen_inst/_0360_ ),
    .B(\wave_gen_inst/_0361_ ),
    .X(\wave_gen_inst/_0362_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3207_  (.A(\wave_gen_inst/_0359_ ),
    .B(\wave_gen_inst/_0362_ ),
    .X(\wave_gen_inst/_0363_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3208_  (.A(\wave_gen_inst/_0343_ ),
    .B(\wave_gen_inst/_0363_ ),
    .X(\wave_gen_inst/_0364_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3209_  (.A(\wave_gen_inst/_0341_ ),
    .B(\wave_gen_inst/_0364_ ),
    .X(\wave_gen_inst/_0365_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3210_  (.A(\wave_gen_inst/_0339_ ),
    .B(\wave_gen_inst/_0365_ ),
    .X(\wave_gen_inst/_0366_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3211_  (.A(\wave_gen_inst/_0338_ ),
    .B(\wave_gen_inst/_0366_ ),
    .Y(\wave_gen_inst/_0367_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3212_  (.A1(\wave_gen_inst/_0337_ ),
    .A2(\wave_gen_inst/_0331_ ),
    .B1(\wave_gen_inst/_0367_ ),
    .Y(\wave_gen_inst/_0368_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3213_  (.A(\wave_gen_inst/_0337_ ),
    .B(\wave_gen_inst/_0331_ ),
    .C(\wave_gen_inst/_0367_ ),
    .Y(\wave_gen_inst/_0369_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3214_  (.A_N(\wave_gen_inst/_0368_ ),
    .B(\wave_gen_inst/_0369_ ),
    .Y(\wave_gen_inst/_0370_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3215_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/_0370_ ),
    .Y(\wave_gen_inst/_0371_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3216_  (.A(\wave_gen_inst/_0336_ ),
    .B(\wave_gen_inst/_0371_ ),
    .Y(\wave_gen_inst/_0372_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3217_  (.A(\wave_gen_inst/_0233_ ),
    .B(\wave_gen_inst/_0372_ ),
    .Y(\wave_gen_inst/_0373_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3219_  (.A(net163),
    .B(\wave_gen_inst/_0111_ ),
    .C(\wave_gen_inst/_0370_ ),
    .X(\wave_gen_inst/_0375_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3220_  (.A1(\wave_gen_inst/param1[5] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[5] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net42),
    .Y(\wave_gen_inst/_0376_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3221_  (.A1(\wave_gen_inst/_0373_ ),
    .A2(\wave_gen_inst/_0375_ ),
    .A3(\wave_gen_inst/_0376_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0004_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3222_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/_0336_ ),
    .C(\wave_gen_inst/_0370_ ),
    .X(\wave_gen_inst/_0377_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3223_  (.A(\wave_gen_inst/_0338_ ),
    .B(\wave_gen_inst/_0366_ ),
    .X(\wave_gen_inst/_0378_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3224_  (.A(\wave_gen_inst/_0378_ ),
    .B(\wave_gen_inst/_0368_ ),
    .Y(\wave_gen_inst/_0379_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3225_  (.A(\wave_gen_inst/_0339_ ),
    .B(\wave_gen_inst/_0365_ ),
    .Y(\wave_gen_inst/_0380_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3226_  (.A(\wave_gen_inst/_0341_ ),
    .B(\wave_gen_inst/_0343_ ),
    .C(\wave_gen_inst/_0363_ ),
    .X(\wave_gen_inst/_0381_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3227_  (.A(\wave_gen_inst/_0345_ ),
    .B(\wave_gen_inst/_0358_ ),
    .C(\wave_gen_inst/_0362_ ),
    .X(\wave_gen_inst/_0382_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3228_  (.A(\wave_gen_inst/_0347_ ),
    .B(\wave_gen_inst/_0346_ ),
    .C(\wave_gen_inst/_0348_ ),
    .X(\wave_gen_inst/_0383_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3229_  (.A_N(\wave_gen_inst/_0351_ ),
    .B(\wave_gen_inst/_0356_ ),
    .Y(\wave_gen_inst/_0384_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3230_  (.A(\wave_gen_inst/_0350_ ),
    .B(\wave_gen_inst/_0357_ ),
    .Y(\wave_gen_inst/_0385_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3231_  (.A(\wave_gen_inst/param1[6] ),
    .B(net480),
    .Y(\wave_gen_inst/_0386_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3232_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0387_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3233_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0388_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3234_  (.A(\wave_gen_inst/_0387_ ),
    .B(\wave_gen_inst/_0388_ ),
    .X(\wave_gen_inst/_0389_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3235_  (.A(\wave_gen_inst/_0386_ ),
    .B(\wave_gen_inst/_0389_ ),
    .Y(\wave_gen_inst/_0390_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3236_  (.A(\wave_gen_inst/_0353_ ),
    .B(\wave_gen_inst/_0352_ ),
    .C(\wave_gen_inst/_0354_ ),
    .X(\wave_gen_inst/_0391_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3237_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0392_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3238_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[6] ),
    .Y(\wave_gen_inst/_0393_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3239_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_0394_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3240_  (.A(\wave_gen_inst/_0393_ ),
    .B(\wave_gen_inst/_0394_ ),
    .X(\wave_gen_inst/_0395_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3241_  (.A(\wave_gen_inst/_0392_ ),
    .B(\wave_gen_inst/_0395_ ),
    .Y(\wave_gen_inst/_0396_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3242_  (.A(\wave_gen_inst/_0391_ ),
    .B(\wave_gen_inst/_0396_ ),
    .Y(\wave_gen_inst/_0397_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3243_  (.A(\wave_gen_inst/_0390_ ),
    .B(\wave_gen_inst/_0397_ ),
    .Y(\wave_gen_inst/_0398_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3244_  (.A(\wave_gen_inst/_0384_ ),
    .B(\wave_gen_inst/_0385_ ),
    .C(\wave_gen_inst/_0398_ ),
    .X(\wave_gen_inst/_0399_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_3245_  (.A1(\wave_gen_inst/_0384_ ),
    .A2(\wave_gen_inst/_0385_ ),
    .B1(\wave_gen_inst/_0398_ ),
    .Y(\wave_gen_inst/_0400_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3246_  (.A(\wave_gen_inst/_0399_ ),
    .B(\wave_gen_inst/_0400_ ),
    .Y(\wave_gen_inst/_0401_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3247_  (.A(\wave_gen_inst/_0383_ ),
    .B(\wave_gen_inst/_0401_ ),
    .Y(\wave_gen_inst/_0402_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3248_  (.A(\wave_gen_inst/_0382_ ),
    .B(\wave_gen_inst/_0402_ ),
    .X(\wave_gen_inst/_0403_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3249_  (.A(\wave_gen_inst/_0250_ ),
    .B(\wave_gen_inst/_0360_ ),
    .Y(\wave_gen_inst/_0404_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3250_  (.A(\wave_gen_inst/param1[5] ),
    .B(net481),
    .C(\wave_gen_inst/_0404_ ),
    .Y(\wave_gen_inst/_0405_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3251_  (.A(\wave_gen_inst/_0405_ ),
    .Y(\wave_gen_inst/_0406_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3252_  (.A(\wave_gen_inst/_0403_ ),
    .B(\wave_gen_inst/_0406_ ),
    .Y(\wave_gen_inst/_0407_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3253_  (.A(\wave_gen_inst/_0381_ ),
    .B(\wave_gen_inst/_0407_ ),
    .X(\wave_gen_inst/_0408_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3254_  (.A(\wave_gen_inst/_0380_ ),
    .B(\wave_gen_inst/_0408_ ),
    .Y(\wave_gen_inst/_0409_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3255_  (.A(\wave_gen_inst/_0379_ ),
    .B(\wave_gen_inst/_0409_ ),
    .Y(\wave_gen_inst/_0410_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3256_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/_0410_ ),
    .Y(\wave_gen_inst/_0411_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3257_  (.A(\wave_gen_inst/_0377_ ),
    .B(\wave_gen_inst/_0411_ ),
    .Y(\wave_gen_inst/_0412_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3258_  (.A(\wave_gen_inst/_0233_ ),
    .B(\wave_gen_inst/_0412_ ),
    .Y(\wave_gen_inst/_0413_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3259_  (.A(net163),
    .B(\wave_gen_inst/_0111_ ),
    .C(\wave_gen_inst/_0410_ ),
    .X(\wave_gen_inst/_0414_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3260_  (.A1(\wave_gen_inst/param1[6] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[6] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net43),
    .Y(\wave_gen_inst/_0415_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3261_  (.A1(\wave_gen_inst/_0413_ ),
    .A2(\wave_gen_inst/_0414_ ),
    .A3(\wave_gen_inst/_0415_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0005_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3262_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/_0377_ ),
    .C(\wave_gen_inst/_0410_ ),
    .X(\wave_gen_inst/_0416_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3263_  (.A(\wave_gen_inst/_0380_ ),
    .B(\wave_gen_inst/_0408_ ),
    .Y(\wave_gen_inst/_0417_ ));
 sky130_fd_sc_hd__o21bai_2 \wave_gen_inst/_3264_  (.A1(\wave_gen_inst/_0378_ ),
    .A2(\wave_gen_inst/_0368_ ),
    .B1_N(\wave_gen_inst/_0409_ ),
    .Y(\wave_gen_inst/_0418_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3265_  (.A(\wave_gen_inst/_0381_ ),
    .B(\wave_gen_inst/_0407_ ),
    .Y(\wave_gen_inst/_0419_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3266_  (.A(\wave_gen_inst/_0382_ ),
    .B(\wave_gen_inst/_0402_ ),
    .Y(\wave_gen_inst/_0420_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3267_  (.A(\wave_gen_inst/_0403_ ),
    .B(\wave_gen_inst/_0406_ ),
    .Y(\wave_gen_inst/_0421_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3268_  (.A(\wave_gen_inst/_0383_ ),
    .B(\wave_gen_inst/_0399_ ),
    .C(\wave_gen_inst/_0400_ ),
    .Y(\wave_gen_inst/_0422_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3269_  (.A(\wave_gen_inst/_0387_ ),
    .B(\wave_gen_inst/_0386_ ),
    .C(\wave_gen_inst/_0388_ ),
    .X(\wave_gen_inst/_0423_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3270_  (.A_N(\wave_gen_inst/_0391_ ),
    .B(\wave_gen_inst/_0396_ ),
    .Y(\wave_gen_inst/_0424_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/_3271_  (.A1(\wave_gen_inst/_0390_ ),
    .A2(\wave_gen_inst/_0397_ ),
    .B1_N(\wave_gen_inst/_0424_ ),
    .Y(\wave_gen_inst/_0425_ ));
 sky130_fd_sc_hd__nand4_2 \wave_gen_inst/_3272_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/param1[8] ),
    .C(\wave_gen_inst/rom_output[10] ),
    .D(net482),
    .Y(\wave_gen_inst/_0426_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3273_  (.A1(\wave_gen_inst/param1[8] ),
    .A2(\wave_gen_inst/rom_output[10] ),
    .B1(net483),
    .B2(\wave_gen_inst/param1[7] ),
    .Y(\wave_gen_inst/_0427_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3274_  (.A(\wave_gen_inst/_0426_ ),
    .SLEEP(\wave_gen_inst/_0427_ ),
    .X(\wave_gen_inst/_0428_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3275_  (.A(\wave_gen_inst/_0393_ ),
    .B(\wave_gen_inst/_0392_ ),
    .C(\wave_gen_inst/_0394_ ),
    .X(\wave_gen_inst/_0429_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3276_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0430_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3277_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[7] ),
    .Y(\wave_gen_inst/_0431_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3278_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0432_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3279_  (.A(\wave_gen_inst/_0431_ ),
    .B(\wave_gen_inst/_0432_ ),
    .X(\wave_gen_inst/_0433_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3280_  (.A(\wave_gen_inst/_0430_ ),
    .B(\wave_gen_inst/_0433_ ),
    .Y(\wave_gen_inst/_0434_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3281_  (.A(\wave_gen_inst/_0429_ ),
    .B(\wave_gen_inst/_0434_ ),
    .Y(\wave_gen_inst/_0435_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3282_  (.A(\wave_gen_inst/_0428_ ),
    .B(\wave_gen_inst/_0435_ ),
    .Y(\wave_gen_inst/_0436_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3283_  (.A(\wave_gen_inst/_0425_ ),
    .B(\wave_gen_inst/_0436_ ),
    .X(\wave_gen_inst/_0437_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3284_  (.A(\wave_gen_inst/_0423_ ),
    .B(\wave_gen_inst/_0437_ ),
    .Y(\wave_gen_inst/_0438_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3285_  (.A1(\wave_gen_inst/_0400_ ),
    .A2(\wave_gen_inst/_0422_ ),
    .B1(\wave_gen_inst/_0438_ ),
    .X(\wave_gen_inst/_0439_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3286_  (.A(\wave_gen_inst/_0400_ ),
    .B(\wave_gen_inst/_0422_ ),
    .C(\wave_gen_inst/_0438_ ),
    .Y(\wave_gen_inst/_0440_ ));
 sky130_fd_sc_hd__or2_0 \wave_gen_inst/_3287_  (.A(\wave_gen_inst/_0439_ ),
    .B(\wave_gen_inst/_0440_ ),
    .X(\wave_gen_inst/_0441_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3288_  (.A1(\wave_gen_inst/_0420_ ),
    .A2(\wave_gen_inst/_0421_ ),
    .B1(\wave_gen_inst/_0441_ ),
    .Y(\wave_gen_inst/_0442_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3289_  (.A(\wave_gen_inst/_0420_ ),
    .B(\wave_gen_inst/_0421_ ),
    .C(\wave_gen_inst/_0441_ ),
    .X(\wave_gen_inst/_0443_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3290_  (.A(\wave_gen_inst/_0442_ ),
    .B(\wave_gen_inst/_0443_ ),
    .Y(\wave_gen_inst/_0444_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3291_  (.A(\wave_gen_inst/_0419_ ),
    .B(\wave_gen_inst/_0444_ ),
    .Y(\wave_gen_inst/_0445_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3292_  (.A1(\wave_gen_inst/_0417_ ),
    .A2(\wave_gen_inst/_0418_ ),
    .B1(\wave_gen_inst/_0445_ ),
    .Y(\wave_gen_inst/_0446_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3293_  (.A(\wave_gen_inst/_0417_ ),
    .B(\wave_gen_inst/_0418_ ),
    .C(\wave_gen_inst/_0445_ ),
    .Y(\wave_gen_inst/_0447_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3294_  (.A_N(\wave_gen_inst/_0446_ ),
    .B(\wave_gen_inst/_0447_ ),
    .Y(\wave_gen_inst/_0448_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3295_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/_0448_ ),
    .Y(\wave_gen_inst/_0449_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3296_  (.A(\wave_gen_inst/_0416_ ),
    .B(\wave_gen_inst/_0449_ ),
    .Y(\wave_gen_inst/_0450_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3300_  (.A1(\wave_gen_inst/param1[7] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(net880),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net44),
    .Y(\wave_gen_inst/_0454_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3301_  (.A1(net163),
    .A2(\wave_gen_inst/_0111_ ),
    .A3(\wave_gen_inst/_0448_ ),
    .B1(\wave_gen_inst/_0454_ ),
    .Y(\wave_gen_inst/_0455_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3302_  (.A1(\wave_gen_inst/_0233_ ),
    .A2(\wave_gen_inst/_0450_ ),
    .B1(\wave_gen_inst/_0455_ ),
    .Y(\wave_gen_inst/_0456_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3303_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0456_ ),
    .Y(\wave_gen_inst/_0006_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3304_  (.A(\wave_gen_inst/_0419_ ),
    .B(\wave_gen_inst/_0444_ ),
    .Y(\wave_gen_inst/_0457_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3305_  (.A(\wave_gen_inst/_0423_ ),
    .B(\wave_gen_inst/_0425_ ),
    .C(\wave_gen_inst/_0436_ ),
    .X(\wave_gen_inst/_0458_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3306_  (.A(\wave_gen_inst/_0434_ ),
    .SLEEP(\wave_gen_inst/_0429_ ),
    .X(\wave_gen_inst/_0459_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3307_  (.A1(\wave_gen_inst/_0428_ ),
    .A2(\wave_gen_inst/_0435_ ),
    .B1(\wave_gen_inst/_0459_ ),
    .Y(\wave_gen_inst/_0460_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3308_  (.A(\wave_gen_inst/param1[8] ),
    .B(net484),
    .Y(\wave_gen_inst/_0461_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3309_  (.A(\wave_gen_inst/_0431_ ),
    .B(\wave_gen_inst/_0430_ ),
    .C(\wave_gen_inst/_0432_ ),
    .X(\wave_gen_inst/_0462_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3310_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0463_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3311_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0464_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3312_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/rom_output[8] ),
    .Y(\wave_gen_inst/_0465_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3313_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[9] ),
    .Y(\wave_gen_inst/_0466_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3314_  (.A(\wave_gen_inst/_0465_ ),
    .B(\wave_gen_inst/_0466_ ),
    .Y(\wave_gen_inst/_0467_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_3315_  (.A1(\wave_gen_inst/_0432_ ),
    .A2(\wave_gen_inst/_0464_ ),
    .B1(\wave_gen_inst/_0467_ ),
    .Y(\wave_gen_inst/_0468_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3316_  (.A(\wave_gen_inst/_0463_ ),
    .B(\wave_gen_inst/_0468_ ),
    .Y(\wave_gen_inst/_0469_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3317_  (.A(\wave_gen_inst/_0462_ ),
    .B(\wave_gen_inst/_0469_ ),
    .Y(\wave_gen_inst/_0470_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3318_  (.A(\wave_gen_inst/_0461_ ),
    .B(\wave_gen_inst/_0470_ ),
    .Y(\wave_gen_inst/_0471_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3319_  (.A(\wave_gen_inst/_0460_ ),
    .B(\wave_gen_inst/_0471_ ),
    .X(\wave_gen_inst/_0472_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3320_  (.A(\wave_gen_inst/_0426_ ),
    .B(\wave_gen_inst/_0472_ ),
    .Y(\wave_gen_inst/_0473_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3321_  (.A(\wave_gen_inst/_0458_ ),
    .B(\wave_gen_inst/_0473_ ),
    .Y(\wave_gen_inst/_0474_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3322_  (.A(\wave_gen_inst/_0442_ ),
    .B(\wave_gen_inst/_0474_ ),
    .X(\wave_gen_inst/_0475_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3323_  (.A(\wave_gen_inst/_0442_ ),
    .B(\wave_gen_inst/_0474_ ),
    .Y(\wave_gen_inst/_0476_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3324_  (.A(\wave_gen_inst/_0475_ ),
    .B(\wave_gen_inst/_0476_ ),
    .Y(\wave_gen_inst/_0477_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3325_  (.A(\wave_gen_inst/_0439_ ),
    .B(\wave_gen_inst/_0477_ ),
    .Y(\wave_gen_inst/_0478_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3326_  (.A1(\wave_gen_inst/_0439_ ),
    .A2(\wave_gen_inst/_0474_ ),
    .B1(\wave_gen_inst/_0478_ ),
    .Y(\wave_gen_inst/_0479_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3327_  (.A(\wave_gen_inst/_0446_ ),
    .B(\wave_gen_inst/_0479_ ),
    .Y(\wave_gen_inst/_0480_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3328_  (.A(\wave_gen_inst/_0479_ ),
    .Y(\wave_gen_inst/_0481_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3329_  (.A(\wave_gen_inst/_0457_ ),
    .B(\wave_gen_inst/_0481_ ),
    .Y(\wave_gen_inst/_0482_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3330_  (.A1(\wave_gen_inst/_0457_ ),
    .A2(\wave_gen_inst/_0480_ ),
    .B1(\wave_gen_inst/_0482_ ),
    .Y(\wave_gen_inst/_0483_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3331_  (.A(\wave_gen_inst/_0112_ ),
    .B(\wave_gen_inst/_0483_ ),
    .Y(\wave_gen_inst/_0484_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3332_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/_0416_ ),
    .C(\wave_gen_inst/_0448_ ),
    .X(\wave_gen_inst/_0485_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3333_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_0483_ ),
    .Y(\wave_gen_inst/_0486_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3334_  (.A(\wave_gen_inst/_0485_ ),
    .B(\wave_gen_inst/_0486_ ),
    .X(\wave_gen_inst/_0487_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3335_  (.A1(\wave_gen_inst/_0485_ ),
    .A2(\wave_gen_inst/_0486_ ),
    .B1(\wave_gen_inst/_0233_ ),
    .Y(\wave_gen_inst/_0488_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3336_  (.A1(\wave_gen_inst/param1[8] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(\wave_gen_inst/counter[8] ),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net45),
    .Y(\wave_gen_inst/_0489_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3337_  (.A1(\wave_gen_inst/_0487_ ),
    .A2(\wave_gen_inst/_0488_ ),
    .B1(\wave_gen_inst/_0489_ ),
    .X(\wave_gen_inst/_0490_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3338_  (.A1(\wave_gen_inst/_0484_ ),
    .A2(\wave_gen_inst/_0490_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0007_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_3339_  (.A1(\wave_gen_inst/_0457_ ),
    .A2(\wave_gen_inst/_0480_ ),
    .B1(\wave_gen_inst/_0482_ ),
    .X(\wave_gen_inst/_0491_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3340_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_0485_ ),
    .C(\wave_gen_inst/_0491_ ),
    .X(\wave_gen_inst/_0492_ ));
 sky130_fd_sc_hd__a211oi_2 \wave_gen_inst/_3341_  (.A1(\wave_gen_inst/_0417_ ),
    .A2(\wave_gen_inst/_0418_ ),
    .B1(\wave_gen_inst/_0445_ ),
    .C1(\wave_gen_inst/_0481_ ),
    .Y(\wave_gen_inst/_0493_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3342_  (.A(\wave_gen_inst/_0475_ ),
    .B(\wave_gen_inst/_0482_ ),
    .C(\wave_gen_inst/_0493_ ),
    .Y(\wave_gen_inst/_0494_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3343_  (.A(\wave_gen_inst/_0473_ ),
    .SLEEP(\wave_gen_inst/_0458_ ),
    .X(\wave_gen_inst/_0495_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3344_  (.A(\wave_gen_inst/_0426_ ),
    .B(\wave_gen_inst/_0460_ ),
    .C(\wave_gen_inst/_0471_ ),
    .X(\wave_gen_inst/_0496_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3345_  (.A(\wave_gen_inst/_0461_ ),
    .B(\wave_gen_inst/_0462_ ),
    .C(\wave_gen_inst/_0469_ ),
    .X(\wave_gen_inst/_0497_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3346_  (.A(\wave_gen_inst/_0465_ ),
    .B(\wave_gen_inst/_0463_ ),
    .C(\wave_gen_inst/_0466_ ),
    .X(\wave_gen_inst/_0498_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3347_  (.A(\wave_gen_inst/param1[9] ),
    .B(net485),
    .Y(\wave_gen_inst/_0499_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3348_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/rom_output[10] ),
    .Y(\wave_gen_inst/_0500_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3349_  (.A(\wave_gen_inst/_0464_ ),
    .B(\wave_gen_inst/_0500_ ),
    .Y(\wave_gen_inst/_0501_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3350_  (.A(\wave_gen_inst/_0499_ ),
    .B(\wave_gen_inst/_0501_ ),
    .Y(\wave_gen_inst/_0502_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3351_  (.A(\wave_gen_inst/_0498_ ),
    .B(\wave_gen_inst/_0502_ ),
    .X(\wave_gen_inst/_0503_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3352_  (.A(\wave_gen_inst/_0497_ ),
    .B(\wave_gen_inst/_0503_ ),
    .Y(\wave_gen_inst/_0504_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3353_  (.A(\wave_gen_inst/_0496_ ),
    .B(\wave_gen_inst/_0504_ ),
    .Y(\wave_gen_inst/_0505_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3354_  (.A(\wave_gen_inst/_0495_ ),
    .B(\wave_gen_inst/_0505_ ),
    .Y(\wave_gen_inst/_0506_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3355_  (.A(\wave_gen_inst/_0495_ ),
    .B(\wave_gen_inst/_0505_ ),
    .X(\wave_gen_inst/_0507_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3356_  (.A(\wave_gen_inst/_0506_ ),
    .B(\wave_gen_inst/_0507_ ),
    .Y(\wave_gen_inst/_0508_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_3357_  (.A1(\wave_gen_inst/_0439_ ),
    .A2(\wave_gen_inst/_0474_ ),
    .B1(\wave_gen_inst/_0508_ ),
    .X(\wave_gen_inst/_0509_ ));
 sky130_fd_sc_hd__nand3_2 \wave_gen_inst/_3358_  (.A(\wave_gen_inst/_0439_ ),
    .B(\wave_gen_inst/_0474_ ),
    .C(\wave_gen_inst/_0508_ ),
    .Y(\wave_gen_inst/_0510_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3359_  (.A(\wave_gen_inst/_0509_ ),
    .B(\wave_gen_inst/_0510_ ),
    .Y(\wave_gen_inst/_0511_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3360_  (.A(\wave_gen_inst/_0494_ ),
    .B(\wave_gen_inst/_0511_ ),
    .Y(\wave_gen_inst/_0512_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3361_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/_0512_ ),
    .X(\wave_gen_inst/_0513_ ));
 sky130_fd_sc_hd__or2_0 \wave_gen_inst/_3362_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/_0512_ ),
    .X(\wave_gen_inst/_0514_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_3363_  (.A(\wave_gen_inst/_0513_ ),
    .B_N(\wave_gen_inst/_0514_ ),
    .Y(\wave_gen_inst/_0515_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3364_  (.A(\wave_gen_inst/_0492_ ),
    .B(\wave_gen_inst/_0515_ ),
    .X(\wave_gen_inst/_0516_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3365_  (.A(\wave_gen_inst/_0233_ ),
    .B(\wave_gen_inst/_0516_ ),
    .Y(\wave_gen_inst/_0517_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3366_  (.A(net163),
    .B(\wave_gen_inst/_0111_ ),
    .C(\wave_gen_inst/_0512_ ),
    .X(\wave_gen_inst/_0518_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3367_  (.A1(\wave_gen_inst/param1[9] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(net829),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net46),
    .Y(\wave_gen_inst/_0519_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3368_  (.A1(\wave_gen_inst/_0517_ ),
    .A2(\wave_gen_inst/_0518_ ),
    .A3(\wave_gen_inst/_0519_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0008_ ));
 sky130_fd_sc_hd__o311ai_2 \wave_gen_inst/_3369_  (.A1(\wave_gen_inst/_0475_ ),
    .A2(\wave_gen_inst/_0482_ ),
    .A3(\wave_gen_inst/_0493_ ),
    .B1(\wave_gen_inst/_0509_ ),
    .C1(\wave_gen_inst/_0510_ ),
    .Y(\wave_gen_inst/_0520_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3370_  (.A(\wave_gen_inst/_0510_ ),
    .B(\wave_gen_inst/_0520_ ),
    .X(\wave_gen_inst/_0521_ ));
 sky130_fd_sc_hd__nand2b_2 \wave_gen_inst/_3371_  (.A_N(\wave_gen_inst/_0496_ ),
    .B(\wave_gen_inst/_0504_ ),
    .Y(\wave_gen_inst/_0522_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3372_  (.A(\wave_gen_inst/_0503_ ),
    .SLEEP(\wave_gen_inst/_0497_ ),
    .X(\wave_gen_inst/_0523_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3373_  (.A(\wave_gen_inst/_0498_ ),
    .B(\wave_gen_inst/_0502_ ),
    .Y(\wave_gen_inst/_0524_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3374_  (.A(\wave_gen_inst/_0464_ ),
    .B(\wave_gen_inst/_0499_ ),
    .C(\wave_gen_inst/_0500_ ),
    .X(\wave_gen_inst/_0525_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3375_  (.A(\wave_gen_inst/param1[11] ),
    .B(net486),
    .Y(\wave_gen_inst/_0526_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3376_  (.A(\wave_gen_inst/_0500_ ),
    .B(\wave_gen_inst/_0526_ ),
    .Y(\wave_gen_inst/_0527_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3377_  (.A1(\wave_gen_inst/param1[11] ),
    .A2(\wave_gen_inst/rom_output[10] ),
    .B1(net487),
    .B2(\wave_gen_inst/param1[10] ),
    .Y(\wave_gen_inst/_0528_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3378_  (.A(\wave_gen_inst/_0525_ ),
    .B(\wave_gen_inst/_0527_ ),
    .C(\wave_gen_inst/_0528_ ),
    .Y(\wave_gen_inst/_0529_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3379_  (.A1(\wave_gen_inst/_0527_ ),
    .A2(\wave_gen_inst/_0528_ ),
    .B1(\wave_gen_inst/_0525_ ),
    .X(\wave_gen_inst/_0530_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3380_  (.A(\wave_gen_inst/_0529_ ),
    .B(\wave_gen_inst/_0530_ ),
    .Y(\wave_gen_inst/_0531_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3381_  (.A(\wave_gen_inst/_0524_ ),
    .B(\wave_gen_inst/_0531_ ),
    .X(\wave_gen_inst/_0532_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3382_  (.A(\wave_gen_inst/_0523_ ),
    .B(\wave_gen_inst/_0532_ ),
    .Y(\wave_gen_inst/_0533_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3383_  (.A(\wave_gen_inst/_0522_ ),
    .B(\wave_gen_inst/_0533_ ),
    .X(\wave_gen_inst/_0534_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3384_  (.A(\wave_gen_inst/_0507_ ),
    .B(\wave_gen_inst/_0534_ ),
    .Y(\wave_gen_inst/_0535_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_3385_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/_0521_ ),
    .C(\wave_gen_inst/_0535_ ),
    .X(\wave_gen_inst/_0536_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3386_  (.A1(\wave_gen_inst/_0513_ ),
    .A2(\wave_gen_inst/_0492_ ),
    .B1(\wave_gen_inst/_0514_ ),
    .Y(\wave_gen_inst/_0537_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3387_  (.A(\wave_gen_inst/_0536_ ),
    .B(\wave_gen_inst/_0537_ ),
    .Y(\wave_gen_inst/_0538_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3388_  (.A(\wave_gen_inst/_0233_ ),
    .B(\wave_gen_inst/_0538_ ),
    .Y(\wave_gen_inst/_0539_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3389_  (.A(\wave_gen_inst/_0521_ ),
    .B(\wave_gen_inst/_0535_ ),
    .Y(\wave_gen_inst/_0540_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3390_  (.A(net163),
    .B(\wave_gen_inst/_0111_ ),
    .C(\wave_gen_inst/_0540_ ),
    .X(\wave_gen_inst/_0541_ ));
 sky130_fd_sc_hd__a222oi_1 \wave_gen_inst/_3391_  (.A1(\wave_gen_inst/param1[10] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0167_ ),
    .B2(net846),
    .C1(\wave_gen_inst/_0169_ ),
    .C2(net16),
    .Y(\wave_gen_inst/_0542_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3392_  (.A1(\wave_gen_inst/_0539_ ),
    .A2(\wave_gen_inst/_0541_ ),
    .A3(\wave_gen_inst/_0542_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0009_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3393_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/_0540_ ),
    .Y(\wave_gen_inst/_0543_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3394_  (.A1(\wave_gen_inst/_0513_ ),
    .A2(\wave_gen_inst/_0492_ ),
    .B1(\wave_gen_inst/_0514_ ),
    .C1(\wave_gen_inst/_0536_ ),
    .Y(\wave_gen_inst/_0544_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3395_  (.A1(\wave_gen_inst/_0510_ ),
    .A2(\wave_gen_inst/_0520_ ),
    .B1(\wave_gen_inst/_0535_ ),
    .Y(\wave_gen_inst/_0545_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_3396_  (.A1(\wave_gen_inst/_0507_ ),
    .A2(\wave_gen_inst/_0534_ ),
    .B1(\wave_gen_inst/_0545_ ),
    .Y(\wave_gen_inst/_0546_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3397_  (.A1(\wave_gen_inst/param1[10] ),
    .A2(\wave_gen_inst/rom_output[10] ),
    .B1(\wave_gen_inst/_0526_ ),
    .Y(\wave_gen_inst/_0547_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3398_  (.A(\wave_gen_inst/_0529_ ),
    .B(\wave_gen_inst/_0547_ ),
    .X(\wave_gen_inst/_0548_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3399_  (.A(\wave_gen_inst/_0524_ ),
    .B(\wave_gen_inst/_0523_ ),
    .C(\wave_gen_inst/_0531_ ),
    .X(\wave_gen_inst/_0549_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3400_  (.A(\wave_gen_inst/_0548_ ),
    .B(\wave_gen_inst/_0549_ ),
    .Y(\wave_gen_inst/_0550_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3401_  (.A(\wave_gen_inst/_0522_ ),
    .B(\wave_gen_inst/_0533_ ),
    .C(\wave_gen_inst/_0550_ ),
    .Y(\wave_gen_inst/_0551_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3402_  (.A1(\wave_gen_inst/_0522_ ),
    .A2(\wave_gen_inst/_0533_ ),
    .B1(\wave_gen_inst/_0550_ ),
    .X(\wave_gen_inst/_0552_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3403_  (.A(\wave_gen_inst/_0551_ ),
    .B(\wave_gen_inst/_0552_ ),
    .Y(\wave_gen_inst/_0553_ ));
 sky130_fd_sc_hd__xnor3_1 \wave_gen_inst/_3404_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_0546_ ),
    .C(\wave_gen_inst/_0553_ ),
    .X(\wave_gen_inst/_0554_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3405_  (.A1(\wave_gen_inst/_0543_ ),
    .A2(\wave_gen_inst/_0544_ ),
    .B1(\wave_gen_inst/_0554_ ),
    .Y(\wave_gen_inst/_0555_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3406_  (.A(\wave_gen_inst/_0543_ ),
    .B(\wave_gen_inst/_0544_ ),
    .C(\wave_gen_inst/_0554_ ),
    .Y(\wave_gen_inst/_0556_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_3407_  (.A_N(\wave_gen_inst/_0555_ ),
    .B(\wave_gen_inst/_0556_ ),
    .C(\wave_gen_inst/_0233_ ),
    .Y(\wave_gen_inst/_0557_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3408_  (.A(\wave_gen_inst/_0546_ ),
    .B(\wave_gen_inst/_0553_ ),
    .X(\wave_gen_inst/_0558_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3409_  (.A(net163),
    .B(\wave_gen_inst/_0111_ ),
    .C(\wave_gen_inst/_0558_ ),
    .X(\wave_gen_inst/_0559_ ));
 sky130_fd_sc_hd__a22o_1 \wave_gen_inst/_3410_  (.A1(\wave_gen_inst/counter[11] ),
    .A2(\wave_gen_inst/_0167_ ),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net17),
    .X(\wave_gen_inst/_0560_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3411_  (.A1(\wave_gen_inst/param1[11] ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/_0560_ ),
    .Y(\wave_gen_inst/_0561_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3412_  (.A1(\wave_gen_inst/_0557_ ),
    .A2(\wave_gen_inst/_0559_ ),
    .A3(\wave_gen_inst/_0561_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0010_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3413_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_0558_ ),
    .X(\wave_gen_inst/_0562_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3414_  (.A(\wave_gen_inst/_0546_ ),
    .B(\wave_gen_inst/_0551_ ),
    .C(\wave_gen_inst/_0552_ ),
    .Y(\wave_gen_inst/_0563_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3415_  (.A(\wave_gen_inst/_0529_ ),
    .B(\wave_gen_inst/_0547_ ),
    .C(\wave_gen_inst/_0549_ ),
    .X(\wave_gen_inst/_0564_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3416_  (.A(\wave_gen_inst/_0527_ ),
    .B(\wave_gen_inst/_0551_ ),
    .C(\wave_gen_inst/_0563_ ),
    .D(\wave_gen_inst/_0564_ ),
    .Y(\wave_gen_inst/_0565_ ));
 sky130_fd_sc_hd__o2111ai_1 \wave_gen_inst/_3417_  (.A1(\wave_gen_inst/_0562_ ),
    .A2(\wave_gen_inst/_0555_ ),
    .B1(\wave_gen_inst/_0565_ ),
    .C1(\wave_gen_inst/_0233_ ),
    .D1(\wave_gen_inst/param1[11] ),
    .Y(\wave_gen_inst/_0566_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3418_  (.A_N(\wave_gen_inst/_0565_ ),
    .B(\wave_gen_inst/_0112_ ),
    .Y(\wave_gen_inst/_0567_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3421_  (.A1(\wave_gen_inst/counter[12] ),
    .A2(\wave_gen_inst/_0167_ ),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net18),
    .Y(\wave_gen_inst/_0570_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3422_  (.A1(\wave_gen_inst/_0566_ ),
    .A2(\wave_gen_inst/_0567_ ),
    .A3(\wave_gen_inst/_0570_ ),
    .B1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0011_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3425_  (.A1(\wave_gen_inst/counter[13] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net19),
    .Y(\wave_gen_inst/_0573_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3426_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0573_ ),
    .Y(\wave_gen_inst/_0012_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3427_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net20),
    .Y(\wave_gen_inst/_0574_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3428_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0574_ ),
    .Y(\wave_gen_inst/_0013_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3429_  (.A1(\wave_gen_inst/counter[15] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net21),
    .Y(\wave_gen_inst/_0575_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3430_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0575_ ),
    .Y(\wave_gen_inst/_0014_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3431_  (.A1(\wave_gen_inst/counter[16] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net22),
    .Y(\wave_gen_inst/_0576_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3432_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0576_ ),
    .Y(\wave_gen_inst/_0015_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3433_  (.A1(\wave_gen_inst/counter[17] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net23),
    .Y(\wave_gen_inst/_0577_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3434_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0577_ ),
    .Y(\wave_gen_inst/_0016_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3435_  (.A1(\wave_gen_inst/counter[18] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net24),
    .Y(\wave_gen_inst/_0578_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3436_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0578_ ),
    .Y(\wave_gen_inst/_0017_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3437_  (.A1(net813),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net25),
    .Y(\wave_gen_inst/_0579_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3438_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0579_ ),
    .Y(\wave_gen_inst/_0018_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3439_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net27),
    .Y(\wave_gen_inst/_0580_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3440_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0580_ ),
    .Y(\wave_gen_inst/_0019_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3442_  (.A1(net814),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net28),
    .Y(\wave_gen_inst/_0582_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3443_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0582_ ),
    .Y(\wave_gen_inst/_0020_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3444_  (.A1(net817),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net29),
    .Y(\wave_gen_inst/_0583_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3445_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0583_ ),
    .Y(\wave_gen_inst/_0021_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3446_  (.A1(\wave_gen_inst/counter[23] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net30),
    .Y(\wave_gen_inst/_0584_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3447_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0584_ ),
    .Y(\wave_gen_inst/_0022_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3448_  (.A1(net882),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net31),
    .Y(\wave_gen_inst/_0585_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3449_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0585_ ),
    .Y(\wave_gen_inst/_0023_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3451_  (.A1(net818),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net32),
    .Y(\wave_gen_inst/_0587_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3452_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0587_ ),
    .Y(\wave_gen_inst/_0024_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3454_  (.A1(\wave_gen_inst/counter[26] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net33),
    .Y(\wave_gen_inst/_0589_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3455_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0589_ ),
    .Y(\wave_gen_inst/_0025_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3457_  (.A1(\wave_gen_inst/counter[27] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net34),
    .Y(\wave_gen_inst/_0591_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3458_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0591_ ),
    .Y(\wave_gen_inst/_0026_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3460_  (.A1(\wave_gen_inst/counter[28] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net35),
    .Y(\wave_gen_inst/_0593_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3461_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0593_ ),
    .Y(\wave_gen_inst/_0027_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3463_  (.A1(\wave_gen_inst/counter[29] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net36),
    .Y(\wave_gen_inst/_0595_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3464_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0595_ ),
    .Y(\wave_gen_inst/_0028_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3466_  (.A1(\wave_gen_inst/counter[30] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net38),
    .Y(\wave_gen_inst/_0597_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3467_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0597_ ),
    .Y(\wave_gen_inst/_0029_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3470_  (.A1(\wave_gen_inst/counter[31] ),
    .A2(net142),
    .B1(\wave_gen_inst/_0169_ ),
    .B2(net39),
    .Y(\wave_gen_inst/_0600_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3471_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0600_ ),
    .Y(\wave_gen_inst/_0030_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \wave_gen_inst/_3472_  (.A(net11),
    .SLEEP(net12),
    .X(\wave_gen_inst/_0601_ ));
 sky130_fd_sc_hd__nor3_4 \wave_gen_inst/_3473_  (.A(net13),
    .B(\wave_gen_inst/_1752_ ),
    .C(\wave_gen_inst/_0601_ ),
    .Y(\wave_gen_inst/_0602_ ));
 sky130_fd_sc_hd__xnor2_4 \wave_gen_inst/_3476_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/counter[1] ),
    .Y(\wave_gen_inst/_0605_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3477_  (.A_N(\wave_gen_inst/counter[0] ),
    .B(\wave_gen_inst/param2[0] ),
    .Y(\wave_gen_inst/_0606_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3478_  (.A(\wave_gen_inst/_0605_ ),
    .B(\wave_gen_inst/_0606_ ),
    .Y(\wave_gen_inst/_0607_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3479_  (.A(\wave_gen_inst/param2[11] ),
    .B(\wave_gen_inst/_0124_ ),
    .Y(\wave_gen_inst/_0608_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3480_  (.A(\wave_gen_inst/_1898_ ),
    .B(\wave_gen_inst/_0124_ ),
    .Y(\wave_gen_inst/_0609_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3481_  (.A(\wave_gen_inst/_1898_ ),
    .B(\wave_gen_inst/_0124_ ),
    .Y(\wave_gen_inst/_0610_ ));
 sky130_fd_sc_hd__nand2b_2 \wave_gen_inst/_3482_  (.A_N(\wave_gen_inst/_0609_ ),
    .B(\wave_gen_inst/_0610_ ),
    .Y(\wave_gen_inst/_0611_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3483_  (.A(\wave_gen_inst/param2[7] ),
    .SLEEP(\wave_gen_inst/counter[7] ),
    .X(\wave_gen_inst/_0612_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3484_  (.A(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/_0141_ ),
    .Y(\wave_gen_inst/_0613_ ));
 sky130_fd_sc_hd__and2_2 \wave_gen_inst/_3485_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/counter[4] ),
    .X(\wave_gen_inst/_0614_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3486_  (.A(\wave_gen_inst/param2[4] ),
    .B(\wave_gen_inst/counter[4] ),
    .Y(\wave_gen_inst/_0615_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_3487_  (.A(\wave_gen_inst/_0614_ ),
    .B(\wave_gen_inst/_0615_ ),
    .Y(\wave_gen_inst/_0616_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3488_  (.A(\wave_gen_inst/_1552_ ),
    .B(\wave_gen_inst/counter[3] ),
    .Y(\wave_gen_inst/_0617_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3489_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/counter[2] ),
    .X(\wave_gen_inst/_0618_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3490_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/counter[2] ),
    .Y(\wave_gen_inst/_0619_ ));
 sky130_fd_sc_hd__or2_2 \wave_gen_inst/_3491_  (.A(\wave_gen_inst/_0618_ ),
    .B(\wave_gen_inst/_0619_ ),
    .X(\wave_gen_inst/_0620_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_3492_  (.A(\wave_gen_inst/_1548_ ),
    .B(\wave_gen_inst/counter[1] ),
    .C(\wave_gen_inst/_0606_ ),
    .X(\wave_gen_inst/_0621_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3493_  (.A(\wave_gen_inst/counter[2] ),
    .SLEEP(\wave_gen_inst/param2[2] ),
    .X(\wave_gen_inst/_0622_ ));
 sky130_fd_sc_hd__a221oi_4 \wave_gen_inst/_3494_  (.A1(\wave_gen_inst/_1552_ ),
    .A2(\wave_gen_inst/counter[3] ),
    .B1(\wave_gen_inst/_0620_ ),
    .B2(\wave_gen_inst/_0621_ ),
    .C1(\wave_gen_inst/_0622_ ),
    .Y(\wave_gen_inst/_0623_ ));
 sky130_fd_sc_hd__o32ai_4 \wave_gen_inst/_3495_  (.A1(\wave_gen_inst/_0616_ ),
    .A2(\wave_gen_inst/_0617_ ),
    .A3(\wave_gen_inst/_0623_ ),
    .B1(\wave_gen_inst/_1578_ ),
    .B2(\wave_gen_inst/param2[4] ),
    .Y(\wave_gen_inst/_0624_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3496_  (.A(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/_0141_ ),
    .Y(\wave_gen_inst/_0625_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_3497_  (.A1(\wave_gen_inst/_0613_ ),
    .A2(\wave_gen_inst/_0624_ ),
    .B1(\wave_gen_inst/_0625_ ),
    .Y(\wave_gen_inst/_0626_ ));
 sky130_fd_sc_hd__maj3_2 \wave_gen_inst/_3498_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/_0135_ ),
    .C(\wave_gen_inst/_0626_ ),
    .X(\wave_gen_inst/_0627_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3499_  (.A_N(\wave_gen_inst/param2[7] ),
    .B(\wave_gen_inst/counter[7] ),
    .Y(\wave_gen_inst/_0628_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_3500_  (.A1(\wave_gen_inst/_0612_ ),
    .A2(\wave_gen_inst/_0627_ ),
    .B1(\wave_gen_inst/_0628_ ),
    .Y(\wave_gen_inst/_0629_ ));
 sky130_fd_sc_hd__xnor2_4 \wave_gen_inst/_3501_  (.A(\wave_gen_inst/param2[9] ),
    .B(\wave_gen_inst/counter[9] ),
    .Y(\wave_gen_inst/_0630_ ));
 sky130_fd_sc_hd__xnor2_4 \wave_gen_inst/_3502_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/counter[8] ),
    .Y(\wave_gen_inst/_0631_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3503_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/_1590_ ),
    .Y(\wave_gen_inst/_0632_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3504_  (.A(\wave_gen_inst/_0630_ ),
    .B(\wave_gen_inst/_0632_ ),
    .Y(\wave_gen_inst/_0633_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_3505_  (.A1(\wave_gen_inst/param2[9] ),
    .A2(\wave_gen_inst/_1646_ ),
    .B1(\wave_gen_inst/_0633_ ),
    .Y(\wave_gen_inst/_0634_ ));
 sky130_fd_sc_hd__a31oi_4 \wave_gen_inst/_3506_  (.A1(\wave_gen_inst/_0629_ ),
    .A2(\wave_gen_inst/_0630_ ),
    .A3(\wave_gen_inst/_0631_ ),
    .B1(\wave_gen_inst/_0634_ ),
    .Y(\wave_gen_inst/_0635_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3507_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/_0123_ ),
    .C(\wave_gen_inst/_0635_ ),
    .X(\wave_gen_inst/_0636_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3508_  (.A(\wave_gen_inst/_0611_ ),
    .SLEEP(\wave_gen_inst/_0636_ ),
    .X(\wave_gen_inst/_0637_ ));
 sky130_fd_sc_hd__or3_2 \wave_gen_inst/_3509_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/_0608_ ),
    .C(\wave_gen_inst/_0637_ ),
    .X(\wave_gen_inst/_0638_ ));
 sky130_fd_sc_hd__or2_4 \wave_gen_inst/_3510_  (.A(\wave_gen_inst/_0149_ ),
    .B(\wave_gen_inst/_0638_ ),
    .X(\wave_gen_inst/_0639_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3512_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_0156_ ),
    .C(\wave_gen_inst/_0639_ ),
    .Y(\wave_gen_inst/_0641_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3513_  (.A(\wave_gen_inst/_0151_ ),
    .B(\wave_gen_inst/_0641_ ),
    .Y(\wave_gen_inst/_0642_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3514_  (.A(\wave_gen_inst/counter[26] ),
    .B(\wave_gen_inst/_0642_ ),
    .Y(\wave_gen_inst/_0643_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3515_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_0643_ ),
    .Y(\wave_gen_inst/_0644_ ));
 sky130_fd_sc_hd__or4_2 \wave_gen_inst/_3516_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/counter[19] ),
    .C(\wave_gen_inst/_0154_ ),
    .D(\wave_gen_inst/_0639_ ),
    .X(\wave_gen_inst/_0645_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3517_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/counter[21] ),
    .C(\wave_gen_inst/_0645_ ),
    .X(\wave_gen_inst/_0646_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3518_  (.A(\wave_gen_inst/_0156_ ),
    .B(\wave_gen_inst/_0639_ ),
    .Y(\wave_gen_inst/_0647_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3519_  (.A1(\wave_gen_inst/counter[22] ),
    .A2(\wave_gen_inst/_0646_ ),
    .B1(\wave_gen_inst/_0647_ ),
    .Y(\wave_gen_inst/_0648_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3520_  (.A1(\wave_gen_inst/counter[16] ),
    .A2(\wave_gen_inst/_0154_ ),
    .A3(\wave_gen_inst/_0639_ ),
    .B1(\wave_gen_inst/counter[19] ),
    .Y(\wave_gen_inst/_0649_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3521_  (.A(\wave_gen_inst/_0649_ ),
    .B(\wave_gen_inst/_0645_ ),
    .X(\wave_gen_inst/_0650_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3522_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_0647_ ),
    .Y(\wave_gen_inst/_0651_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_3523_  (.A_N(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/_0650_ ),
    .C(\wave_gen_inst/_0651_ ),
    .Y(\wave_gen_inst/_0652_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3524_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/_0645_ ),
    .X(\wave_gen_inst/_0653_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3525_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_0639_ ),
    .X(\wave_gen_inst/_0654_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3526_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/_0641_ ),
    .Y(\wave_gen_inst/_0655_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3527_  (.A(\wave_gen_inst/counter[21] ),
    .B(\wave_gen_inst/counter[26] ),
    .C(\wave_gen_inst/counter[29] ),
    .D(\wave_gen_inst/_0154_ ),
    .Y(\wave_gen_inst/_0656_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_3528_  (.A(\wave_gen_inst/_0653_ ),
    .B(\wave_gen_inst/_0654_ ),
    .C(\wave_gen_inst/_0655_ ),
    .D(\wave_gen_inst/_0656_ ),
    .Y(\wave_gen_inst/_0657_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3529_  (.A(\wave_gen_inst/_0652_ ),
    .B(\wave_gen_inst/_0657_ ),
    .Y(\wave_gen_inst/_0658_ ));
 sky130_fd_sc_hd__nand3_2 \wave_gen_inst/_3530_  (.A(\wave_gen_inst/_0644_ ),
    .B(\wave_gen_inst/_0648_ ),
    .C(\wave_gen_inst/_0658_ ),
    .Y(\wave_gen_inst/_0659_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_3531_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/counter[24] ),
    .C(\wave_gen_inst/_0156_ ),
    .D(\wave_gen_inst/_0639_ ),
    .X(\wave_gen_inst/_0660_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3532_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/counter[26] ),
    .C(\wave_gen_inst/counter[27] ),
    .D(\wave_gen_inst/_0660_ ),
    .Y(\wave_gen_inst/_0661_ ));
 sky130_fd_sc_hd__nand2b_2 \wave_gen_inst/_3533_  (.A_N(\wave_gen_inst/counter[28] ),
    .B(\wave_gen_inst/_0661_ ),
    .Y(\wave_gen_inst/_0662_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3534_  (.A_N(\wave_gen_inst/_0661_ ),
    .B(\wave_gen_inst/counter[28] ),
    .Y(\wave_gen_inst/_0663_ ));
 sky130_fd_sc_hd__nand4bb_2 \wave_gen_inst/_3535_  (.A_N(\wave_gen_inst/counter[30] ),
    .B_N(\wave_gen_inst/counter[31] ),
    .C(\wave_gen_inst/_0662_ ),
    .D(\wave_gen_inst/_0663_ ),
    .Y(\wave_gen_inst/_0664_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3536_  (.A(\wave_gen_inst/_0659_ ),
    .B(\wave_gen_inst/_0664_ ),
    .Y(\wave_gen_inst/_0665_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3537_  (.A(\wave_gen_inst/counter[0] ),
    .B(\wave_gen_inst/counter[1] ),
    .Y(\wave_gen_inst/_0666_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3538_  (.A(\wave_gen_inst/counter[6] ),
    .B(\wave_gen_inst/counter[7] ),
    .C(\wave_gen_inst/counter[8] ),
    .D(\wave_gen_inst/counter[11] ),
    .Y(\wave_gen_inst/_0667_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_3539_  (.A(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/counter[3] ),
    .C(\wave_gen_inst/counter[4] ),
    .D(\wave_gen_inst/counter[5] ),
    .X(\wave_gen_inst/_0668_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3540_  (.A(\wave_gen_inst/counter[9] ),
    .B(\wave_gen_inst/counter[10] ),
    .C(\wave_gen_inst/_0668_ ),
    .Y(\wave_gen_inst/_0669_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3541_  (.A(\wave_gen_inst/_0161_ ),
    .B(\wave_gen_inst/_0667_ ),
    .C(\wave_gen_inst/_0669_ ),
    .X(\wave_gen_inst/_0670_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3542_  (.A(\wave_gen_inst/_0666_ ),
    .B(\wave_gen_inst/_0670_ ),
    .Y(\wave_gen_inst/_0671_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3543_  (.A(\wave_gen_inst/_0611_ ),
    .B(\wave_gen_inst/_0636_ ),
    .X(\wave_gen_inst/_0672_ ));
 sky130_fd_sc_hd__xor2_4 \wave_gen_inst/_3544_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/counter[10] ),
    .X(\wave_gen_inst/_0673_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3545_  (.A(\wave_gen_inst/_0673_ ),
    .B(\wave_gen_inst/_0635_ ),
    .Y(\wave_gen_inst/_0674_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3546_  (.A(\wave_gen_inst/param2[9] ),
    .B(\wave_gen_inst/counter[9] ),
    .Y(\wave_gen_inst/_0675_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3547_  (.A(\wave_gen_inst/param2[9] ),
    .B(\wave_gen_inst/counter[9] ),
    .Y(\wave_gen_inst/_0676_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \wave_gen_inst/_3548_  (.A(\wave_gen_inst/_0675_ ),
    .SLEEP(\wave_gen_inst/_0676_ ),
    .X(\wave_gen_inst/_0677_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3549_  (.A1(\wave_gen_inst/_0629_ ),
    .A2(\wave_gen_inst/_0631_ ),
    .B1(\wave_gen_inst/_0632_ ),
    .Y(\wave_gen_inst/_0678_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3550_  (.A(\wave_gen_inst/_0677_ ),
    .B(\wave_gen_inst/_0678_ ),
    .Y(\wave_gen_inst/_0679_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3551_  (.A(\wave_gen_inst/_0629_ ),
    .B(\wave_gen_inst/_0631_ ),
    .Y(\wave_gen_inst/_0680_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3552_  (.A(\wave_gen_inst/param2[7] ),
    .B(\wave_gen_inst/counter[7] ),
    .Y(\wave_gen_inst/_0681_ ));
 sky130_fd_sc_hd__or2_1 \wave_gen_inst/_3553_  (.A(\wave_gen_inst/param2[7] ),
    .B(\wave_gen_inst/counter[7] ),
    .X(\wave_gen_inst/_0682_ ));
 sky130_fd_sc_hd__and2_2 \wave_gen_inst/_3554_  (.A(\wave_gen_inst/_0681_ ),
    .B(\wave_gen_inst/_0682_ ),
    .X(\wave_gen_inst/_0683_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3556_  (.A(\wave_gen_inst/_0627_ ),
    .B(\wave_gen_inst/_0683_ ),
    .Y(\wave_gen_inst/_0685_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3557_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/counter[6] ),
    .X(\wave_gen_inst/_0686_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3558_  (.A(\wave_gen_inst/_0686_ ),
    .B(\wave_gen_inst/_0626_ ),
    .Y(\wave_gen_inst/_0687_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3559_  (.A(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/counter[5] ),
    .X(\wave_gen_inst/_0688_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_3560_  (.A(\wave_gen_inst/param2[5] ),
    .B(\wave_gen_inst/counter[5] ),
    .Y(\wave_gen_inst/_0689_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_3561_  (.A(\wave_gen_inst/_0688_ ),
    .B(\wave_gen_inst/_0689_ ),
    .Y(\wave_gen_inst/_0690_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3562_  (.A(\wave_gen_inst/_0624_ ),
    .B(\wave_gen_inst/_0690_ ),
    .X(\wave_gen_inst/_0691_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3563_  (.A(\wave_gen_inst/_0617_ ),
    .B(\wave_gen_inst/_0623_ ),
    .Y(\wave_gen_inst/_0692_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3564_  (.A(\wave_gen_inst/_0616_ ),
    .B(\wave_gen_inst/_0692_ ),
    .X(\wave_gen_inst/_0693_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3565_  (.A1(\wave_gen_inst/_0620_ ),
    .A2(\wave_gen_inst/_0621_ ),
    .B1(\wave_gen_inst/_0622_ ),
    .Y(\wave_gen_inst/_0694_ ));
 sky130_fd_sc_hd__xor2_4 \wave_gen_inst/_3566_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/counter[3] ),
    .X(\wave_gen_inst/_0695_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3567_  (.A(\wave_gen_inst/_0694_ ),
    .B(\wave_gen_inst/_0695_ ),
    .Y(\wave_gen_inst/_0696_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3568_  (.A(\wave_gen_inst/_0620_ ),
    .B(\wave_gen_inst/_0621_ ),
    .Y(\wave_gen_inst/_0697_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3569_  (.A(\wave_gen_inst/_0607_ ),
    .Y(\wave_gen_inst/_0698_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3570_  (.A(\wave_gen_inst/_1672_ ),
    .B(\wave_gen_inst/_0606_ ),
    .X(\wave_gen_inst/_0699_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3571_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/param1[1] ),
    .C(\wave_gen_inst/_0699_ ),
    .Y(\wave_gen_inst/_0700_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3572_  (.A1(\wave_gen_inst/param1[0] ),
    .A2(\wave_gen_inst/_0699_ ),
    .B1(\wave_gen_inst/param1[1] ),
    .Y(\wave_gen_inst/_0701_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3573_  (.A1(\wave_gen_inst/_0698_ ),
    .A2(\wave_gen_inst/_0700_ ),
    .B1(\wave_gen_inst/_0701_ ),
    .Y(\wave_gen_inst/_0702_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3574_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/_0697_ ),
    .C(\wave_gen_inst/_0702_ ),
    .X(\wave_gen_inst/_0703_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3575_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/_0696_ ),
    .C(\wave_gen_inst/_0703_ ),
    .X(\wave_gen_inst/_0704_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3576_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/_0693_ ),
    .C(\wave_gen_inst/_0704_ ),
    .X(\wave_gen_inst/_0705_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3577_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/_0691_ ),
    .C(\wave_gen_inst/_0705_ ),
    .X(\wave_gen_inst/_0706_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3578_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/_0687_ ),
    .C(\wave_gen_inst/_0706_ ),
    .X(\wave_gen_inst/_0707_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3579_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_0685_ ),
    .C(\wave_gen_inst/_0707_ ),
    .X(\wave_gen_inst/_0708_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3580_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/_0680_ ),
    .C(\wave_gen_inst/_0708_ ),
    .X(\wave_gen_inst/_0709_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3581_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/_0679_ ),
    .C(\wave_gen_inst/_0709_ ),
    .X(\wave_gen_inst/_0710_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3582_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_0674_ ),
    .C(\wave_gen_inst/_0710_ ),
    .X(\wave_gen_inst/_0711_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3583_  (.A1(\wave_gen_inst/param1[11] ),
    .A2(\wave_gen_inst/_0672_ ),
    .B1(\wave_gen_inst/_0711_ ),
    .Y(\wave_gen_inst/_0712_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3584_  (.A1(\wave_gen_inst/_0608_ ),
    .A2(\wave_gen_inst/_0637_ ),
    .B1(\wave_gen_inst/counter[12] ),
    .Y(\wave_gen_inst/_0713_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3585_  (.A(\wave_gen_inst/_0638_ ),
    .B(\wave_gen_inst/_0713_ ),
    .X(\wave_gen_inst/_0714_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_3586_  (.A(\wave_gen_inst/_0149_ ),
    .B_N(\wave_gen_inst/_0714_ ),
    .Y(\wave_gen_inst/_0715_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3587_  (.A1(\wave_gen_inst/param1[11] ),
    .A2(\wave_gen_inst/_0672_ ),
    .B1(\wave_gen_inst/_0715_ ),
    .Y(\wave_gen_inst/_0716_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3588_  (.A(\wave_gen_inst/_0712_ ),
    .B(\wave_gen_inst/_0716_ ),
    .Y(\wave_gen_inst/_0717_ ));
 sky130_fd_sc_hd__and3_4 \wave_gen_inst/_3589_  (.A(\wave_gen_inst/_0665_ ),
    .B(\wave_gen_inst/_0671_ ),
    .C(\wave_gen_inst/_0717_ ),
    .X(\wave_gen_inst/_0718_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3591_  (.A1(\wave_gen_inst/param1[1] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_0720_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3592_  (.A1(\wave_gen_inst/_0607_ ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_0720_ ),
    .Y(\wave_gen_inst/_0721_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_3593_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/counter[8] ),
    .X(\wave_gen_inst/_0722_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_3594_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/counter[6] ),
    .Y(\wave_gen_inst/_0723_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3595_  (.A(\wave_gen_inst/_1552_ ),
    .B(\wave_gen_inst/_1655_ ),
    .Y(\wave_gen_inst/_0724_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_3596_  (.A(\wave_gen_inst/_0618_ ),
    .B(\wave_gen_inst/_0619_ ),
    .Y(\wave_gen_inst/_0725_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3597_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_0726_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3598_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/counter[1] ),
    .Y(\wave_gen_inst/_0727_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_3599_  (.A1(\wave_gen_inst/_0605_ ),
    .A2(\wave_gen_inst/_0726_ ),
    .B1(\wave_gen_inst/_0727_ ),
    .Y(\wave_gen_inst/_0728_ ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/_3600_  (.A1(\wave_gen_inst/param2[3] ),
    .A2(\wave_gen_inst/counter[3] ),
    .B1(\wave_gen_inst/_0725_ ),
    .B2(\wave_gen_inst/_0728_ ),
    .C1(\wave_gen_inst/_0618_ ),
    .X(\wave_gen_inst/_0729_ ));
 sky130_fd_sc_hd__a311oi_4 \wave_gen_inst/_3601_  (.A1(\wave_gen_inst/_0616_ ),
    .A2(\wave_gen_inst/_0724_ ),
    .A3(\wave_gen_inst/_0729_ ),
    .B1(\wave_gen_inst/_0688_ ),
    .C1(\wave_gen_inst/_0614_ ),
    .Y(\wave_gen_inst/_0730_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3602_  (.A(\wave_gen_inst/param2[6] ),
    .B(\wave_gen_inst/counter[6] ),
    .Y(\wave_gen_inst/_0731_ ));
 sky130_fd_sc_hd__o311ai_4 \wave_gen_inst/_3603_  (.A1(\wave_gen_inst/_0723_ ),
    .A2(\wave_gen_inst/_0689_ ),
    .A3(\wave_gen_inst/_0730_ ),
    .B1(\wave_gen_inst/_0681_ ),
    .C1(\wave_gen_inst/_0731_ ),
    .Y(\wave_gen_inst/_0732_ ));
 sky130_fd_sc_hd__a32oi_4 \wave_gen_inst/_3604_  (.A1(\wave_gen_inst/_0722_ ),
    .A2(\wave_gen_inst/_0682_ ),
    .A3(\wave_gen_inst/_0732_ ),
    .B1(\wave_gen_inst/counter[8] ),
    .B2(\wave_gen_inst/param2[8] ),
    .Y(\wave_gen_inst/_0733_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3605_  (.A1(\wave_gen_inst/_0675_ ),
    .A2(\wave_gen_inst/_0733_ ),
    .B1(\wave_gen_inst/_0676_ ),
    .Y(\wave_gen_inst/_0734_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3606_  (.A(\wave_gen_inst/param2[10] ),
    .B(net968),
    .C(\wave_gen_inst/_0734_ ),
    .X(\wave_gen_inst/_0735_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_3607_  (.A1(\wave_gen_inst/_0609_ ),
    .A2(\wave_gen_inst/_0735_ ),
    .B1(\wave_gen_inst/_0610_ ),
    .Y(\wave_gen_inst/_0736_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3608_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/counter[13] ),
    .C(\wave_gen_inst/counter[14] ),
    .X(\wave_gen_inst/_0737_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_3609_  (.A(\wave_gen_inst/counter[15] ),
    .B(\wave_gen_inst/_0737_ ),
    .Y(\wave_gen_inst/_0738_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3610_  (.A(\wave_gen_inst/_0736_ ),
    .B(\wave_gen_inst/_0738_ ),
    .Y(\wave_gen_inst/_0739_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3611_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/counter[17] ),
    .C(\wave_gen_inst/counter[18] ),
    .X(\wave_gen_inst/_0740_ ));
 sky130_fd_sc_hd__and3_2 \wave_gen_inst/_3612_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_0739_ ),
    .C(\wave_gen_inst/_0740_ ),
    .X(\wave_gen_inst/_0741_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3614_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/counter[21] ),
    .C(\wave_gen_inst/_0741_ ),
    .X(\wave_gen_inst/_0743_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3615_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/counter[23] ),
    .C(\wave_gen_inst/_0743_ ),
    .Y(\wave_gen_inst/_0744_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3616_  (.A(\wave_gen_inst/counter[24] ),
    .SLEEP(\wave_gen_inst/_0744_ ),
    .X(\wave_gen_inst/_0745_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3617_  (.A1(\wave_gen_inst/counter[25] ),
    .A2(\wave_gen_inst/_0745_ ),
    .B1(\wave_gen_inst/counter[26] ),
    .Y(\wave_gen_inst/_0746_ ));
 sky130_fd_sc_hd__and3_2 \wave_gen_inst/_3618_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/counter[21] ),
    .C(\wave_gen_inst/counter[22] ),
    .X(\wave_gen_inst/_0747_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3619_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/counter[25] ),
    .C(\wave_gen_inst/counter[26] ),
    .X(\wave_gen_inst/_0748_ ));
 sky130_fd_sc_hd__and4_1 \wave_gen_inst/_3620_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_0747_ ),
    .C(\wave_gen_inst/_0741_ ),
    .D(\wave_gen_inst/_0748_ ),
    .X(\wave_gen_inst/_0749_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3621_  (.A(\wave_gen_inst/_0746_ ),
    .B(\wave_gen_inst/_0749_ ),
    .Y(\wave_gen_inst/_0750_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3622_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/_0743_ ),
    .Y(\wave_gen_inst/_0751_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_3623_  (.A1(\wave_gen_inst/_0747_ ),
    .A2(\wave_gen_inst/_0741_ ),
    .B1(\wave_gen_inst/_0751_ ),
    .Y(\wave_gen_inst/_0752_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3624_  (.A(\wave_gen_inst/counter[28] ),
    .B(\wave_gen_inst/counter[29] ),
    .Y(\wave_gen_inst/_0753_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_3625_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/counter[26] ),
    .C(\wave_gen_inst/counter[27] ),
    .D(\wave_gen_inst/_0745_ ),
    .Y(\wave_gen_inst/_0754_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3626_  (.A(\wave_gen_inst/_0753_ ),
    .B(\wave_gen_inst/_0754_ ),
    .Y(\wave_gen_inst/_0755_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3627_  (.A1(\wave_gen_inst/counter[30] ),
    .A2(\wave_gen_inst/_0755_ ),
    .B1(\wave_gen_inst/counter[31] ),
    .Y(\wave_gen_inst/_0756_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3628_  (.A1(\wave_gen_inst/counter[30] ),
    .A2(\wave_gen_inst/counter[31] ),
    .A3(\wave_gen_inst/_0755_ ),
    .B1(\wave_gen_inst/_0756_ ),
    .Y(\wave_gen_inst/_0757_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3629_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_0749_ ),
    .Y(\wave_gen_inst/_0758_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3630_  (.A_N(\wave_gen_inst/_0757_ ),
    .B(\wave_gen_inst/_0758_ ),
    .Y(\wave_gen_inst/_0759_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_3631_  (.A(\wave_gen_inst/counter[17] ),
    .B(\wave_gen_inst/counter[18] ),
    .Y(\wave_gen_inst/_0760_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3632_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_0739_ ),
    .Y(\wave_gen_inst/_0761_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3633_  (.A(\wave_gen_inst/_0760_ ),
    .B(\wave_gen_inst/_0761_ ),
    .Y(\wave_gen_inst/_0762_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3634_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_0762_ ),
    .Y(\wave_gen_inst/_0763_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3635_  (.A(\wave_gen_inst/_0741_ ),
    .B(\wave_gen_inst/_0763_ ),
    .Y(\wave_gen_inst/_0764_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3636_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_0739_ ),
    .X(\wave_gen_inst/_0765_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3637_  (.A_N(\wave_gen_inst/_0736_ ),
    .B(\wave_gen_inst/counter[12] ),
    .Y(\wave_gen_inst/_0766_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3638_  (.A(\wave_gen_inst/counter[13] ),
    .SLEEP(\wave_gen_inst/_0766_ ),
    .X(\wave_gen_inst/_0767_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3639_  (.A(\wave_gen_inst/counter[14] ),
    .B(\wave_gen_inst/_0767_ ),
    .Y(\wave_gen_inst/_0768_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3640_  (.A(\wave_gen_inst/counter[15] ),
    .B(\wave_gen_inst/_0768_ ),
    .Y(\wave_gen_inst/_0769_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3641_  (.A(\wave_gen_inst/counter[14] ),
    .B(\wave_gen_inst/_0767_ ),
    .Y(\wave_gen_inst/_0770_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3642_  (.A(\wave_gen_inst/counter[13] ),
    .B(\wave_gen_inst/_0766_ ),
    .X(\wave_gen_inst/_0771_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3643_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/_0736_ ),
    .X(\wave_gen_inst/_0772_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3644_  (.A(\wave_gen_inst/_0611_ ),
    .B(\wave_gen_inst/_0735_ ),
    .X(\wave_gen_inst/_0773_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3645_  (.A(\wave_gen_inst/_0673_ ),
    .B(\wave_gen_inst/_0734_ ),
    .Y(\wave_gen_inst/_0774_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3646_  (.A(\wave_gen_inst/_0630_ ),
    .B(\wave_gen_inst/_0733_ ),
    .Y(\wave_gen_inst/_0775_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3647_  (.A(\wave_gen_inst/_0682_ ),
    .B(\wave_gen_inst/_0732_ ),
    .X(\wave_gen_inst/_0776_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3648_  (.A(\wave_gen_inst/_0722_ ),
    .B(\wave_gen_inst/_0776_ ),
    .Y(\wave_gen_inst/_0777_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3649_  (.A(\wave_gen_inst/_0723_ ),
    .B(\wave_gen_inst/_0689_ ),
    .C(\wave_gen_inst/_0730_ ),
    .X(\wave_gen_inst/_0778_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3650_  (.A(\wave_gen_inst/_0731_ ),
    .B(\wave_gen_inst/_0778_ ),
    .Y(\wave_gen_inst/_0779_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3651_  (.A(\wave_gen_inst/_0683_ ),
    .B(\wave_gen_inst/_0779_ ),
    .Y(\wave_gen_inst/_0780_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3652_  (.A1(\wave_gen_inst/_0689_ ),
    .A2(\wave_gen_inst/_0730_ ),
    .B1(\wave_gen_inst/_0723_ ),
    .Y(\wave_gen_inst/_0781_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3653_  (.A(\wave_gen_inst/_0778_ ),
    .B(\wave_gen_inst/_0781_ ),
    .Y(\wave_gen_inst/_0782_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3654_  (.A(\wave_gen_inst/_0724_ ),
    .B(\wave_gen_inst/_0729_ ),
    .X(\wave_gen_inst/_0783_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_3655_  (.A1(\wave_gen_inst/_0616_ ),
    .A2(\wave_gen_inst/_0783_ ),
    .B1(\wave_gen_inst/_0614_ ),
    .X(\wave_gen_inst/_0784_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3656_  (.A(\wave_gen_inst/_0690_ ),
    .B(\wave_gen_inst/_0784_ ),
    .Y(\wave_gen_inst/_0785_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3657_  (.A(\wave_gen_inst/_0616_ ),
    .B(\wave_gen_inst/_0783_ ),
    .Y(\wave_gen_inst/_0786_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_3658_  (.A1(\wave_gen_inst/_0725_ ),
    .A2(\wave_gen_inst/_0728_ ),
    .B1(\wave_gen_inst/_0618_ ),
    .X(\wave_gen_inst/_0787_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3659_  (.A(\wave_gen_inst/_0695_ ),
    .B(\wave_gen_inst/_0787_ ),
    .Y(\wave_gen_inst/_0788_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3660_  (.A(\wave_gen_inst/_0605_ ),
    .B(\wave_gen_inst/_0726_ ),
    .X(\wave_gen_inst/_0789_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3661_  (.A1(\wave_gen_inst/_0700_ ),
    .A2(\wave_gen_inst/_0789_ ),
    .B1(\wave_gen_inst/_0701_ ),
    .Y(\wave_gen_inst/_0790_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3662_  (.A(\wave_gen_inst/_0725_ ),
    .B(\wave_gen_inst/_0728_ ),
    .Y(\wave_gen_inst/_0791_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3663_  (.A(\wave_gen_inst/param1[2] ),
    .B(\wave_gen_inst/_0790_ ),
    .C(\wave_gen_inst/_0791_ ),
    .X(\wave_gen_inst/_0792_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3664_  (.A(\wave_gen_inst/param1[3] ),
    .B(\wave_gen_inst/_0788_ ),
    .C(\wave_gen_inst/_0792_ ),
    .X(\wave_gen_inst/_0793_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3665_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/_0786_ ),
    .C(\wave_gen_inst/_0793_ ),
    .X(\wave_gen_inst/_0794_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3666_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/_0785_ ),
    .C(\wave_gen_inst/_0794_ ),
    .X(\wave_gen_inst/_0795_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3667_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/_0782_ ),
    .C(\wave_gen_inst/_0795_ ),
    .X(\wave_gen_inst/_0796_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3668_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_0780_ ),
    .C(\wave_gen_inst/_0796_ ),
    .X(\wave_gen_inst/_0797_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3669_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/_0777_ ),
    .C(\wave_gen_inst/_0797_ ),
    .X(\wave_gen_inst/_0798_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3670_  (.A(\wave_gen_inst/param1[9] ),
    .B(\wave_gen_inst/_0775_ ),
    .C(\wave_gen_inst/_0798_ ),
    .X(\wave_gen_inst/_0799_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3671_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_0774_ ),
    .C(\wave_gen_inst/_0799_ ),
    .X(\wave_gen_inst/_0800_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3672_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/_0773_ ),
    .C(\wave_gen_inst/_0800_ ),
    .X(\wave_gen_inst/_0801_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_3673_  (.A(\wave_gen_inst/_0770_ ),
    .B(\wave_gen_inst/_0771_ ),
    .C(\wave_gen_inst/_0772_ ),
    .D(\wave_gen_inst/_0801_ ),
    .Y(\wave_gen_inst/_0802_ ));
 sky130_fd_sc_hd__or4_1 \wave_gen_inst/_3674_  (.A(\wave_gen_inst/_0764_ ),
    .B(\wave_gen_inst/_0765_ ),
    .C(\wave_gen_inst/_0769_ ),
    .D(\wave_gen_inst/_0802_ ),
    .X(\wave_gen_inst/_0803_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3675_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/_0745_ ),
    .X(\wave_gen_inst/_0804_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3676_  (.A1(\wave_gen_inst/_0747_ ),
    .A2(\wave_gen_inst/_0741_ ),
    .B1(\wave_gen_inst/counter[23] ),
    .Y(\wave_gen_inst/_0805_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3677_  (.A(\wave_gen_inst/_0744_ ),
    .SLEEP(\wave_gen_inst/_0805_ ),
    .X(\wave_gen_inst/_0806_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3678_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/counter[28] ),
    .C(\wave_gen_inst/_0749_ ),
    .Y(\wave_gen_inst/_0807_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3679_  (.A(\wave_gen_inst/counter[29] ),
    .B(\wave_gen_inst/_0807_ ),
    .X(\wave_gen_inst/_0808_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3680_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/_0744_ ),
    .X(\wave_gen_inst/_0809_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3681_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/_0741_ ),
    .Y(\wave_gen_inst/_0810_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3682_  (.A(\wave_gen_inst/counter[17] ),
    .B(\wave_gen_inst/_0761_ ),
    .X(\wave_gen_inst/_0811_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_3683_  (.A(\wave_gen_inst/_0808_ ),
    .B(\wave_gen_inst/_0809_ ),
    .C(\wave_gen_inst/_0810_ ),
    .D(\wave_gen_inst/_0811_ ),
    .Y(\wave_gen_inst/_0812_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3684_  (.A(\wave_gen_inst/_0803_ ),
    .B(\wave_gen_inst/_0804_ ),
    .C(\wave_gen_inst/_0806_ ),
    .D(\wave_gen_inst/_0812_ ),
    .Y(\wave_gen_inst/_0813_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3685_  (.A(\wave_gen_inst/counter[30] ),
    .B(\wave_gen_inst/_0755_ ),
    .Y(\wave_gen_inst/_0814_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3686_  (.A(\wave_gen_inst/counter[28] ),
    .B(\wave_gen_inst/_0754_ ),
    .Y(\wave_gen_inst/_0815_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3687_  (.A1(\wave_gen_inst/counter[16] ),
    .A2(\wave_gen_inst/counter[17] ),
    .A3(\wave_gen_inst/_0739_ ),
    .B1(\wave_gen_inst/counter[18] ),
    .Y(\wave_gen_inst/_0816_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3688_  (.A(\wave_gen_inst/_0762_ ),
    .B(\wave_gen_inst/_0816_ ),
    .Y(\wave_gen_inst/_0817_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3689_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(\wave_gen_inst/_0741_ ),
    .B1(\wave_gen_inst/counter[21] ),
    .Y(\wave_gen_inst/_0818_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3690_  (.A(\wave_gen_inst/_0743_ ),
    .B(\wave_gen_inst/_0818_ ),
    .Y(\wave_gen_inst/_0819_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3691_  (.A(\wave_gen_inst/_0815_ ),
    .B(\wave_gen_inst/_0817_ ),
    .C(\wave_gen_inst/_0819_ ),
    .Y(\wave_gen_inst/_0820_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3692_  (.A(\wave_gen_inst/_0813_ ),
    .B(\wave_gen_inst/_0814_ ),
    .C(\wave_gen_inst/_0820_ ),
    .Y(\wave_gen_inst/_0821_ ));
 sky130_fd_sc_hd__or4_4 \wave_gen_inst/_3693_  (.A(\wave_gen_inst/_0750_ ),
    .B(\wave_gen_inst/_0752_ ),
    .C(\wave_gen_inst/_0759_ ),
    .D(\wave_gen_inst/_0821_ ),
    .X(\wave_gen_inst/_0822_ ));
 sky130_fd_sc_hd__nor3b_1 \wave_gen_inst/_3696_  (.A(\wave_gen_inst/_0822_ ),
    .B(\wave_gen_inst/sign ),
    .C_N(\wave_gen_inst/_0789_ ),
    .Y(\wave_gen_inst/_0825_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3697_  (.A1(\wave_gen_inst/_0721_ ),
    .A2(\wave_gen_inst/_0825_ ),
    .B1(\wave_gen_inst/_1753_ ),
    .Y(\wave_gen_inst/_0826_ ));
 sky130_fd_sc_hd__nand2_8 \wave_gen_inst/_3700_  (.A(net13),
    .B(\wave_gen_inst/_0601_ ),
    .Y(\wave_gen_inst/_0829_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3702_  (.A1(net163),
    .A2(\wave_gen_inst/_0607_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_0831_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3703_  (.A1(net163),
    .A2(\wave_gen_inst/_0789_ ),
    .B1(\wave_gen_inst/_0831_ ),
    .Y(\wave_gen_inst/_0832_ ));
 sky130_fd_sc_hd__or3_4 \wave_gen_inst/_3704_  (.A(net13),
    .B(\wave_gen_inst/_1752_ ),
    .C(\wave_gen_inst/_0601_ ),
    .X(\wave_gen_inst/_0833_ ));
 sky130_fd_sc_hd__o2111a_1 \wave_gen_inst/_3707_  (.A1(\wave_gen_inst/counter[1] ),
    .A2(\wave_gen_inst/_0111_ ),
    .B1(\wave_gen_inst/_0826_ ),
    .C1(\wave_gen_inst/_0832_ ),
    .D1(\wave_gen_inst/_0833_ ),
    .X(\wave_gen_inst/_0836_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3708_  (.A(\wave_gen_inst/_1663_ ),
    .B(\wave_gen_inst/_1705_ ),
    .Y(\wave_gen_inst/_0837_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3709_  (.A(\wave_gen_inst/_1555_ ),
    .B(\wave_gen_inst/_0837_ ),
    .Y(\wave_gen_inst/_0838_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3710_  (.A1(\wave_gen_inst/_1526_ ),
    .A2(\wave_gen_inst/_0838_ ),
    .B1(\wave_gen_inst/_0161_ ),
    .Y(\wave_gen_inst/_0839_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3711_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/param2[4] ),
    .C(\wave_gen_inst/_0837_ ),
    .Y(\wave_gen_inst/_0840_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3712_  (.A(\wave_gen_inst/_0690_ ),
    .B(\wave_gen_inst/_0840_ ),
    .X(\wave_gen_inst/_0841_ ));
 sky130_fd_sc_hd__nand4_4 \wave_gen_inst/_3713_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/counter[23] ),
    .C(\wave_gen_inst/_0747_ ),
    .D(\wave_gen_inst/_0740_ ),
    .Y(\wave_gen_inst/_0842_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3714_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_0748_ ),
    .Y(\wave_gen_inst/_0843_ ));
 sky130_fd_sc_hd__nand4_2 \wave_gen_inst/_3715_  (.A(\wave_gen_inst/counter[28] ),
    .B(\wave_gen_inst/counter[29] ),
    .C(\wave_gen_inst/counter[30] ),
    .D(\wave_gen_inst/counter[31] ),
    .Y(\wave_gen_inst/_0844_ ));
 sky130_fd_sc_hd__nor4_4 \wave_gen_inst/_3716_  (.A(\wave_gen_inst/_0738_ ),
    .B(\wave_gen_inst/_0842_ ),
    .C(\wave_gen_inst/_0843_ ),
    .D(\wave_gen_inst/_0844_ ),
    .Y(\wave_gen_inst/_0845_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_3717_  (.A(\wave_gen_inst/_1526_ ),
    .B(\wave_gen_inst/_0838_ ),
    .Y(\wave_gen_inst/_0846_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_3718_  (.A(\wave_gen_inst/_0605_ ),
    .B(\wave_gen_inst/_0606_ ),
    .X(\wave_gen_inst/_0847_ ));
 sky130_fd_sc_hd__nor3_2 \wave_gen_inst/_3719_  (.A(\wave_gen_inst/param2[0] ),
    .B(\wave_gen_inst/param2[1] ),
    .C(\wave_gen_inst/param2[2] ),
    .Y(\wave_gen_inst/_0848_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3720_  (.A(\wave_gen_inst/_0695_ ),
    .B(\wave_gen_inst/_0848_ ),
    .Y(\wave_gen_inst/_0849_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3721_  (.A(\wave_gen_inst/_1723_ ),
    .B(\wave_gen_inst/_0848_ ),
    .Y(\wave_gen_inst/_0850_ ));
 sky130_fd_sc_hd__o32ai_1 \wave_gen_inst/_3722_  (.A1(\wave_gen_inst/param2[6] ),
    .A2(\wave_gen_inst/param2[7] ),
    .A3(\wave_gen_inst/_0850_ ),
    .B1(\wave_gen_inst/_0722_ ),
    .B2(\wave_gen_inst/_0677_ ),
    .Y(\wave_gen_inst/_0851_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3723_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_0837_ ),
    .Y(\wave_gen_inst/_0852_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3724_  (.A(\wave_gen_inst/_0616_ ),
    .B(\wave_gen_inst/_0852_ ),
    .Y(\wave_gen_inst/_0853_ ));
 sky130_fd_sc_hd__o221ai_1 \wave_gen_inst/_3725_  (.A1(\wave_gen_inst/_1525_ ),
    .A2(\wave_gen_inst/_0673_ ),
    .B1(\wave_gen_inst/_0683_ ),
    .B2(\wave_gen_inst/param2[6] ),
    .C1(\wave_gen_inst/_0686_ ),
    .Y(\wave_gen_inst/_0854_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_3726_  (.A1(\wave_gen_inst/param2[6] ),
    .A2(\wave_gen_inst/_0683_ ),
    .B1(\wave_gen_inst/_0838_ ),
    .B2(\wave_gen_inst/_0854_ ),
    .Y(\wave_gen_inst/_0855_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_3727_  (.A(\wave_gen_inst/_0849_ ),
    .B(\wave_gen_inst/_0851_ ),
    .C(\wave_gen_inst/_0853_ ),
    .D(\wave_gen_inst/_0855_ ),
    .Y(\wave_gen_inst/_0856_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3728_  (.A(\wave_gen_inst/param2[8] ),
    .B(\wave_gen_inst/counter[8] ),
    .Y(\wave_gen_inst/_0857_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3729_  (.A1(\wave_gen_inst/counter[8] ),
    .A2(\wave_gen_inst/_0630_ ),
    .B1(\wave_gen_inst/_0857_ ),
    .Y(\wave_gen_inst/_0858_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3730_  (.A(\wave_gen_inst/_1705_ ),
    .B(\wave_gen_inst/_0725_ ),
    .Y(\wave_gen_inst/_0859_ ));
 sky130_fd_sc_hd__o41ai_1 \wave_gen_inst/_3731_  (.A1(\wave_gen_inst/param2[6] ),
    .A2(\wave_gen_inst/param2[7] ),
    .A3(\wave_gen_inst/_0850_ ),
    .A4(\wave_gen_inst/_0858_ ),
    .B1(\wave_gen_inst/_0859_ ),
    .Y(\wave_gen_inst/_0860_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3732_  (.A(\wave_gen_inst/_0686_ ),
    .B(\wave_gen_inst/_0683_ ),
    .Y(\wave_gen_inst/_0861_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3733_  (.A1(\wave_gen_inst/_1531_ ),
    .A2(\wave_gen_inst/counter[0] ),
    .B1(\wave_gen_inst/_0605_ ),
    .Y(\wave_gen_inst/_0862_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3734_  (.A1(\wave_gen_inst/param2[8] ),
    .A2(\wave_gen_inst/_0677_ ),
    .B1(\wave_gen_inst/_0862_ ),
    .Y(\wave_gen_inst/_0863_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3735_  (.A1(\wave_gen_inst/_0838_ ),
    .A2(\wave_gen_inst/_0861_ ),
    .B1(\wave_gen_inst/_0863_ ),
    .Y(\wave_gen_inst/_0864_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3736_  (.A(\wave_gen_inst/_0847_ ),
    .B(\wave_gen_inst/_0856_ ),
    .C(\wave_gen_inst/_0860_ ),
    .D(\wave_gen_inst/_0864_ ),
    .Y(\wave_gen_inst/_0865_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3737_  (.A(\wave_gen_inst/param2[10] ),
    .B(\wave_gen_inst/_1525_ ),
    .C(\wave_gen_inst/_0850_ ),
    .Y(\wave_gen_inst/_0866_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3738_  (.A(\wave_gen_inst/_0611_ ),
    .B(\wave_gen_inst/_0866_ ),
    .X(\wave_gen_inst/_0867_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3739_  (.A1(\wave_gen_inst/_1525_ ),
    .A2(\wave_gen_inst/_0850_ ),
    .B1(\wave_gen_inst/_0673_ ),
    .Y(\wave_gen_inst/_0868_ ));
 sky130_fd_sc_hd__o2111ai_1 \wave_gen_inst/_3740_  (.A1(\wave_gen_inst/_0845_ ),
    .A2(\wave_gen_inst/_0846_ ),
    .B1(\wave_gen_inst/_0865_ ),
    .C1(\wave_gen_inst/_0867_ ),
    .D1(\wave_gen_inst/_0868_ ),
    .Y(\wave_gen_inst/_0869_ ));
 sky130_fd_sc_hd__or3_2 \wave_gen_inst/_3741_  (.A(\wave_gen_inst/_0839_ ),
    .B(\wave_gen_inst/_0841_ ),
    .C(\wave_gen_inst/_0869_ ),
    .X(\wave_gen_inst/_0870_ ));
 sky130_fd_sc_hd__nand4_4 \wave_gen_inst/_3742_  (.A(\wave_gen_inst/_1901_ ),
    .B(\wave_gen_inst/_1814_ ),
    .C(\wave_gen_inst/_1816_ ),
    .D(\wave_gen_inst/_1818_ ),
    .Y(\wave_gen_inst/_0871_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3743_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/param1[5] ),
    .C(\wave_gen_inst/param1[6] ),
    .D(\wave_gen_inst/_0871_ ),
    .Y(\wave_gen_inst/_0872_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3744_  (.A_N(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_0872_ ),
    .Y(\wave_gen_inst/_0873_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3745_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/param1[9] ),
    .C(\wave_gen_inst/_0873_ ),
    .Y(\wave_gen_inst/_0874_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_3746_  (.A_N(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_0874_ ),
    .Y(\wave_gen_inst/_0875_ ));
 sky130_fd_sc_hd__or2_1 \wave_gen_inst/_3747_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/_0875_ ),
    .X(\wave_gen_inst/_0876_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3748_  (.A(\wave_gen_inst/param1[11] ),
    .B(\wave_gen_inst/_0875_ ),
    .Y(\wave_gen_inst/_0877_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3749_  (.A(\wave_gen_inst/counter[11] ),
    .B(\wave_gen_inst/_0877_ ),
    .Y(\wave_gen_inst/_0878_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3750_  (.A(\wave_gen_inst/_0161_ ),
    .B(\wave_gen_inst/_0878_ ),
    .Y(\wave_gen_inst/_0879_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3751_  (.A1(\wave_gen_inst/param1[8] ),
    .A2(\wave_gen_inst/_0873_ ),
    .B1(\wave_gen_inst/param1[9] ),
    .X(\wave_gen_inst/_0880_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3752_  (.A(\wave_gen_inst/_0874_ ),
    .B(\wave_gen_inst/_0880_ ),
    .Y(\wave_gen_inst/_0881_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3753_  (.A(\wave_gen_inst/_1646_ ),
    .B(\wave_gen_inst/_0881_ ),
    .Y(\wave_gen_inst/_0882_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3754_  (.A(\wave_gen_inst/param1[10] ),
    .B(\wave_gen_inst/_0874_ ),
    .Y(\wave_gen_inst/_0883_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3755_  (.A(\wave_gen_inst/_0123_ ),
    .B(\wave_gen_inst/_0883_ ),
    .Y(\wave_gen_inst/_0884_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3756_  (.A1(\wave_gen_inst/_0876_ ),
    .A2(\wave_gen_inst/_0877_ ),
    .B1(\wave_gen_inst/counter[11] ),
    .Y(\wave_gen_inst/_0885_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3757_  (.A(\wave_gen_inst/_0876_ ),
    .B(\wave_gen_inst/_0845_ ),
    .Y(\wave_gen_inst/_0886_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3758_  (.A(\wave_gen_inst/param1[8] ),
    .B(\wave_gen_inst/_0873_ ),
    .X(\wave_gen_inst/_0887_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3759_  (.A(\wave_gen_inst/counter[8] ),
    .B(\wave_gen_inst/_0887_ ),
    .Y(\wave_gen_inst/_0888_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3760_  (.A(\wave_gen_inst/param1[7] ),
    .B(\wave_gen_inst/_0872_ ),
    .Y(\wave_gen_inst/_0889_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3761_  (.A(\wave_gen_inst/_0133_ ),
    .B(\wave_gen_inst/_0889_ ),
    .Y(\wave_gen_inst/_0890_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3762_  (.A(\wave_gen_inst/_0888_ ),
    .B(\wave_gen_inst/_0890_ ),
    .Y(\wave_gen_inst/_0891_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3763_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/param1[5] ),
    .C(\wave_gen_inst/_0871_ ),
    .Y(\wave_gen_inst/_0892_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3764_  (.A(\wave_gen_inst/param1[6] ),
    .B(\wave_gen_inst/_0892_ ),
    .Y(\wave_gen_inst/_0893_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3765_  (.A(\wave_gen_inst/_0135_ ),
    .B(\wave_gen_inst/_0893_ ),
    .Y(\wave_gen_inst/_0894_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3766_  (.A(\wave_gen_inst/param1[1] ),
    .B(\wave_gen_inst/counter[1] ),
    .Y(\wave_gen_inst/_0895_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3767_  (.A(\wave_gen_inst/_1901_ ),
    .B(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_0896_ ));
 sky130_fd_sc_hd__nor3b_1 \wave_gen_inst/_3768_  (.A(\wave_gen_inst/_0895_ ),
    .B(\wave_gen_inst/param1[0] ),
    .C_N(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_0897_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3769_  (.A1(\wave_gen_inst/_0895_ ),
    .A2(\wave_gen_inst/_0896_ ),
    .B1(\wave_gen_inst/_0897_ ),
    .Y(\wave_gen_inst/_0898_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3770_  (.A(\wave_gen_inst/_1901_ ),
    .B(\wave_gen_inst/_1814_ ),
    .C(\wave_gen_inst/_1816_ ),
    .Y(\wave_gen_inst/_0899_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3771_  (.A1(\wave_gen_inst/param1[0] ),
    .A2(\wave_gen_inst/param1[1] ),
    .B1(\wave_gen_inst/param1[2] ),
    .Y(\wave_gen_inst/_0900_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3772_  (.A(\wave_gen_inst/_0899_ ),
    .B(\wave_gen_inst/_0900_ ),
    .Y(\wave_gen_inst/_0901_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3773_  (.A(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/_0901_ ),
    .X(\wave_gen_inst/_0902_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3774_  (.A(\wave_gen_inst/_1818_ ),
    .B(\wave_gen_inst/_0899_ ),
    .Y(\wave_gen_inst/_0903_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3775_  (.A(\wave_gen_inst/counter[3] ),
    .B(\wave_gen_inst/_0903_ ),
    .Y(\wave_gen_inst/_0904_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3776_  (.A(\wave_gen_inst/param1[4] ),
    .B(\wave_gen_inst/_0871_ ),
    .X(\wave_gen_inst/_0905_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3777_  (.A(\wave_gen_inst/counter[4] ),
    .B(\wave_gen_inst/_0905_ ),
    .Y(\wave_gen_inst/_0906_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3778_  (.A(\wave_gen_inst/_0898_ ),
    .B(\wave_gen_inst/_0902_ ),
    .C(\wave_gen_inst/_0904_ ),
    .D(\wave_gen_inst/_0906_ ),
    .Y(\wave_gen_inst/_0907_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_3779_  (.A1(\wave_gen_inst/param1[4] ),
    .A2(\wave_gen_inst/_0871_ ),
    .B1(\wave_gen_inst/param1[5] ),
    .X(\wave_gen_inst/_0908_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3780_  (.A(\wave_gen_inst/_0892_ ),
    .B(\wave_gen_inst/_0908_ ),
    .Y(\wave_gen_inst/_0909_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3781_  (.A(\wave_gen_inst/_0141_ ),
    .B(\wave_gen_inst/_0909_ ),
    .Y(\wave_gen_inst/_0910_ ));
 sky130_fd_sc_hd__o2111ai_2 \wave_gen_inst/_3782_  (.A1(\wave_gen_inst/counter[8] ),
    .A2(\wave_gen_inst/_0887_ ),
    .B1(\wave_gen_inst/_0894_ ),
    .C1(\wave_gen_inst/_0907_ ),
    .D1(\wave_gen_inst/_0910_ ),
    .Y(\wave_gen_inst/_0911_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3783_  (.A(\wave_gen_inst/_0885_ ),
    .B(\wave_gen_inst/_0886_ ),
    .C(\wave_gen_inst/_0891_ ),
    .D(\wave_gen_inst/_0911_ ),
    .Y(\wave_gen_inst/_0912_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3784_  (.A(\wave_gen_inst/_0882_ ),
    .B(\wave_gen_inst/_0884_ ),
    .C(\wave_gen_inst/_0912_ ),
    .Y(\wave_gen_inst/_0913_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_3785_  (.A1(\wave_gen_inst/_0876_ ),
    .A2(\wave_gen_inst/_0879_ ),
    .B1(\wave_gen_inst/_0913_ ),
    .Y(\wave_gen_inst/_0914_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3786_  (.A1(net15),
    .A2(\wave_gen_inst/_0914_ ),
    .B1(\wave_gen_inst/_1833_ ),
    .Y(\wave_gen_inst/_0915_ ));
 sky130_fd_sc_hd__o21a_2 \wave_gen_inst/_3787_  (.A1(net15),
    .A2(\wave_gen_inst/_0870_ ),
    .B1(\wave_gen_inst/_0915_ ),
    .X(\wave_gen_inst/_0916_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3788_  (.A(net13),
    .B(\wave_gen_inst/_0162_ ),
    .C(\wave_gen_inst/_0870_ ),
    .Y(\wave_gen_inst/_0917_ ));
 sky130_fd_sc_hd__o31ai_4 \wave_gen_inst/_3789_  (.A1(net13),
    .A2(\wave_gen_inst/_1752_ ),
    .A3(\wave_gen_inst/_0914_ ),
    .B1(\wave_gen_inst/_0917_ ),
    .Y(\wave_gen_inst/_0918_ ));
 sky130_fd_sc_hd__nor2_8 \wave_gen_inst/_3790_  (.A(\wave_gen_inst/_0916_ ),
    .B(\wave_gen_inst/_0918_ ),
    .Y(\wave_gen_inst/_0919_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3791_  (.A(\wave_gen_inst/counter[0] ),
    .B(net843),
    .Y(\wave_gen_inst/_0920_ ));
 sky130_fd_sc_hd__or3b_1 \wave_gen_inst/_3792_  (.A(\wave_gen_inst/_0666_ ),
    .B(\wave_gen_inst/_0919_ ),
    .C_N(\wave_gen_inst/_0920_ ),
    .X(\wave_gen_inst/_0921_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/_3793_  (.A1(\wave_gen_inst/_1671_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_0836_ ),
    .B2(\wave_gen_inst/_0921_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0031_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3797_  (.A(\wave_gen_inst/_0697_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_0925_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3798_  (.A1(\wave_gen_inst/param1[2] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_0925_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_0926_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3799_  (.A1(\wave_gen_inst/sign ),
    .A2(\wave_gen_inst/_0791_ ),
    .A3(\wave_gen_inst/_0822_ ),
    .B1(\wave_gen_inst/_0926_ ),
    .Y(\wave_gen_inst/_0927_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3801_  (.A(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/_0920_ ),
    .X(\wave_gen_inst/_0929_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3802_  (.A(\wave_gen_inst/counter[2] ),
    .B(net163),
    .X(\wave_gen_inst/_0930_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3803_  (.A1(\wave_gen_inst/counter[1] ),
    .A2(\wave_gen_inst/_0930_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_0931_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3804_  (.A1(\wave_gen_inst/counter[1] ),
    .A2(\wave_gen_inst/_0930_ ),
    .B1(\wave_gen_inst/_0931_ ),
    .Y(\wave_gen_inst/_0932_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3806_  (.A(\wave_gen_inst/_0232_ ),
    .B(\wave_gen_inst/_0791_ ),
    .Y(\wave_gen_inst/_0934_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3807_  (.A1(net163),
    .A2(\wave_gen_inst/_0697_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_0935_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3808_  (.A1(\wave_gen_inst/_0934_ ),
    .A2(\wave_gen_inst/_0935_ ),
    .B1(net141),
    .Y(\wave_gen_inst/_0936_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3809_  (.A1(\wave_gen_inst/_0919_ ),
    .A2(\wave_gen_inst/_0929_ ),
    .B1(\wave_gen_inst/_0932_ ),
    .C1(\wave_gen_inst/_0936_ ),
    .Y(\wave_gen_inst/_0937_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3810_  (.A1(\wave_gen_inst/_1753_ ),
    .A2(\wave_gen_inst/_0927_ ),
    .B1(\wave_gen_inst/_0937_ ),
    .Y(\wave_gen_inst/_0938_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3812_  (.A(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_0940_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3813_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_0938_ ),
    .C(\wave_gen_inst/_0940_ ),
    .Y(\wave_gen_inst/_0032_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3814_  (.A(\wave_gen_inst/_0696_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_0941_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3815_  (.A1(\wave_gen_inst/param1[3] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_0941_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_0942_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3816_  (.A(\wave_gen_inst/sign ),
    .B(\wave_gen_inst/_0788_ ),
    .C(\wave_gen_inst/_0822_ ),
    .X(\wave_gen_inst/_0943_ ));
 sky130_fd_sc_hd__nand2_4 \wave_gen_inst/_3817_  (.A(net13),
    .B(\wave_gen_inst/_1752_ ),
    .Y(\wave_gen_inst/_0944_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3818_  (.A1(\wave_gen_inst/_0942_ ),
    .A2(\wave_gen_inst/_0943_ ),
    .B1(\wave_gen_inst/_0944_ ),
    .Y(\wave_gen_inst/_0945_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3819_  (.A1(\wave_gen_inst/counter[0] ),
    .A2(\wave_gen_inst/counter[1] ),
    .A3(\wave_gen_inst/counter[2] ),
    .B1(\wave_gen_inst/counter[3] ),
    .Y(\wave_gen_inst/_0946_ ));
 sky130_fd_sc_hd__nand4_2 \wave_gen_inst/_3820_  (.A(\wave_gen_inst/counter[0] ),
    .B(\wave_gen_inst/counter[1] ),
    .C(\wave_gen_inst/counter[2] ),
    .D(\wave_gen_inst/counter[3] ),
    .Y(\wave_gen_inst/_0947_ ));
 sky130_fd_sc_hd__nor3b_1 \wave_gen_inst/_3821_  (.A(\wave_gen_inst/_0919_ ),
    .B(\wave_gen_inst/_0946_ ),
    .C_N(\wave_gen_inst/_0947_ ),
    .Y(\wave_gen_inst/_0948_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3823_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0788_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_0950_ ));
 sky130_fd_sc_hd__a21boi_0 \wave_gen_inst/_3824_  (.A1(net163),
    .A2(\wave_gen_inst/_0696_ ),
    .B1_N(\wave_gen_inst/_0950_ ),
    .Y(\wave_gen_inst/_0951_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_3825_  (.A(\wave_gen_inst/counter[1] ),
    .B(\wave_gen_inst/counter[2] ),
    .C(net163),
    .X(\wave_gen_inst/_0952_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3826_  (.A(\wave_gen_inst/counter[3] ),
    .B(net163),
    .X(\wave_gen_inst/_0953_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3827_  (.A(\wave_gen_inst/_0952_ ),
    .B(\wave_gen_inst/_0953_ ),
    .X(\wave_gen_inst/_0954_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3828_  (.A1(\wave_gen_inst/_0952_ ),
    .A2(\wave_gen_inst/_0953_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_0955_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3829_  (.A1(\wave_gen_inst/_0954_ ),
    .A2(\wave_gen_inst/_0955_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_0956_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3830_  (.A(\wave_gen_inst/_0945_ ),
    .B(\wave_gen_inst/_0948_ ),
    .C(\wave_gen_inst/_0951_ ),
    .D(\wave_gen_inst/_0956_ ),
    .Y(\wave_gen_inst/_0957_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3831_  (.A1(\wave_gen_inst/_1655_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_0957_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0033_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3832_  (.A(\wave_gen_inst/_0693_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_0958_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3833_  (.A1(\wave_gen_inst/param1[4] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_0958_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_0959_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3834_  (.A1(\wave_gen_inst/sign ),
    .A2(\wave_gen_inst/_0786_ ),
    .A3(\wave_gen_inst/_0822_ ),
    .B1(\wave_gen_inst/_0959_ ),
    .Y(\wave_gen_inst/_0960_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3835_  (.A(\wave_gen_inst/_1578_ ),
    .B(\wave_gen_inst/_0947_ ),
    .Y(\wave_gen_inst/_0961_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3837_  (.A(\wave_gen_inst/counter[3] ),
    .B(net163),
    .X(\wave_gen_inst/_0963_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3838_  (.A(\wave_gen_inst/_0963_ ),
    .B(\wave_gen_inst/_0954_ ),
    .Y(\wave_gen_inst/_0964_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3839_  (.A(\wave_gen_inst/counter[4] ),
    .B(net163),
    .X(\wave_gen_inst/_0965_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3840_  (.A(\wave_gen_inst/counter[4] ),
    .B(net163),
    .Y(\wave_gen_inst/_0966_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3841_  (.A(\wave_gen_inst/_0964_ ),
    .B(\wave_gen_inst/_0965_ ),
    .C(\wave_gen_inst/_0966_ ),
    .X(\wave_gen_inst/_0967_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3842_  (.A1(\wave_gen_inst/_0965_ ),
    .A2(\wave_gen_inst/_0966_ ),
    .B1(\wave_gen_inst/_0964_ ),
    .Y(\wave_gen_inst/_0968_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_3843_  (.A(net13),
    .B(net11),
    .Y(\wave_gen_inst/_0969_ ));
 sky130_fd_sc_hd__nor2_4 \wave_gen_inst/_3844_  (.A(net12),
    .B(\wave_gen_inst/_0969_ ),
    .Y(\wave_gen_inst/_0970_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3845_  (.A(\wave_gen_inst/_0232_ ),
    .B(\wave_gen_inst/_0786_ ),
    .Y(\wave_gen_inst/_0971_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3846_  (.A(\wave_gen_inst/_0970_ ),
    .B(\wave_gen_inst/_0971_ ),
    .Y(\wave_gen_inst/_0972_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3847_  (.A1(net163),
    .A2(\wave_gen_inst/_0693_ ),
    .B1(\wave_gen_inst/_0972_ ),
    .Y(\wave_gen_inst/_0973_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_3848_  (.A1(\wave_gen_inst/_0106_ ),
    .A2(\wave_gen_inst/_0967_ ),
    .A3(\wave_gen_inst/_0968_ ),
    .B1(net141),
    .C1(\wave_gen_inst/_0973_ ),
    .Y(\wave_gen_inst/_0974_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3849_  (.A1(\wave_gen_inst/_0919_ ),
    .A2(\wave_gen_inst/_0961_ ),
    .B1(\wave_gen_inst/_0974_ ),
    .Y(\wave_gen_inst/_0975_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3850_  (.A1(\wave_gen_inst/_1753_ ),
    .A2(\wave_gen_inst/_0960_ ),
    .B1(\wave_gen_inst/_0975_ ),
    .Y(\wave_gen_inst/_0976_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3851_  (.A1(\wave_gen_inst/_1578_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_0976_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0034_ ));
 sky130_fd_sc_hd__or2_0 \wave_gen_inst/_3852_  (.A(\wave_gen_inst/param1[5] ),
    .B(\wave_gen_inst/_0718_ ),
    .X(\wave_gen_inst/_0977_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3853_  (.A(\wave_gen_inst/_0691_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_0978_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3854_  (.A(\wave_gen_inst/sign ),
    .B(\wave_gen_inst/_0785_ ),
    .C(\wave_gen_inst/_0822_ ),
    .Y(\wave_gen_inst/_0979_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3855_  (.A1(\wave_gen_inst/sign ),
    .A2(\wave_gen_inst/_0977_ ),
    .A3(\wave_gen_inst/_0978_ ),
    .B1(\wave_gen_inst/_0979_ ),
    .Y(\wave_gen_inst/_0980_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3856_  (.A(\wave_gen_inst/_1578_ ),
    .B(\wave_gen_inst/_0947_ ),
    .Y(\wave_gen_inst/_0981_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3857_  (.A(\wave_gen_inst/counter[5] ),
    .B(\wave_gen_inst/_0981_ ),
    .Y(\wave_gen_inst/_0982_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3858_  (.A(net163),
    .B(\wave_gen_inst/_0691_ ),
    .Y(\wave_gen_inst/_0983_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3859_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0785_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_0984_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3860_  (.A(\wave_gen_inst/counter[5] ),
    .B(net163),
    .Y(\wave_gen_inst/_0985_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3861_  (.A(\wave_gen_inst/counter[5] ),
    .B(net163),
    .Y(\wave_gen_inst/_0986_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_3862_  (.A(\wave_gen_inst/_0985_ ),
    .SLEEP(\wave_gen_inst/_0986_ ),
    .X(\wave_gen_inst/_0987_ ));
 sky130_fd_sc_hd__a211oi_2 \wave_gen_inst/_3863_  (.A1(\wave_gen_inst/_0952_ ),
    .A2(\wave_gen_inst/_0953_ ),
    .B1(\wave_gen_inst/_0965_ ),
    .C1(\wave_gen_inst/_0963_ ),
    .Y(\wave_gen_inst/_0988_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3864_  (.A(\wave_gen_inst/_0966_ ),
    .B(\wave_gen_inst/_0988_ ),
    .Y(\wave_gen_inst/_0989_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3865_  (.A1(\wave_gen_inst/_0987_ ),
    .A2(\wave_gen_inst/_0989_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_0990_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3866_  (.A1(\wave_gen_inst/_0987_ ),
    .A2(\wave_gen_inst/_0989_ ),
    .B1(\wave_gen_inst/_0990_ ),
    .Y(\wave_gen_inst/_0991_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3867_  (.A1(\wave_gen_inst/_0983_ ),
    .A2(\wave_gen_inst/_0984_ ),
    .B1(\wave_gen_inst/_0991_ ),
    .C1(net141),
    .Y(\wave_gen_inst/_0992_ ));
 sky130_fd_sc_hd__o221a_1 \wave_gen_inst/_3868_  (.A1(\wave_gen_inst/_0944_ ),
    .A2(\wave_gen_inst/_0980_ ),
    .B1(\wave_gen_inst/_0982_ ),
    .B2(\wave_gen_inst/_0919_ ),
    .C1(\wave_gen_inst/_0992_ ),
    .X(\wave_gen_inst/_0993_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3869_  (.A1(\wave_gen_inst/_0141_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_0993_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0035_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3870_  (.A(\wave_gen_inst/_0687_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_0994_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3871_  (.A1(\wave_gen_inst/param1[6] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_0994_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_0995_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3872_  (.A1(\wave_gen_inst/sign ),
    .A2(\wave_gen_inst/_0782_ ),
    .A3(\wave_gen_inst/_0822_ ),
    .B1(\wave_gen_inst/_0995_ ),
    .Y(\wave_gen_inst/_0996_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3873_  (.A(\wave_gen_inst/_1753_ ),
    .B(\wave_gen_inst/_0996_ ),
    .Y(\wave_gen_inst/_0997_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3874_  (.A(\wave_gen_inst/counter[5] ),
    .B(\wave_gen_inst/_0981_ ),
    .Y(\wave_gen_inst/_0998_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3875_  (.A(\wave_gen_inst/_0135_ ),
    .B(\wave_gen_inst/_0998_ ),
    .Y(\wave_gen_inst/_0999_ ));
 sky130_fd_sc_hd__nand3_2 \wave_gen_inst/_3876_  (.A(\wave_gen_inst/counter[5] ),
    .B(\wave_gen_inst/counter[6] ),
    .C(\wave_gen_inst/_0981_ ),
    .Y(\wave_gen_inst/_1000_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3877_  (.A(\wave_gen_inst/_0999_ ),
    .B(\wave_gen_inst/_1000_ ),
    .Y(\wave_gen_inst/_1001_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3878_  (.A(\wave_gen_inst/_0919_ ),
    .B(\wave_gen_inst/_1001_ ),
    .Y(\wave_gen_inst/_1002_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3879_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0782_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1003_ ));
 sky130_fd_sc_hd__a21boi_0 \wave_gen_inst/_3880_  (.A1(net163),
    .A2(\wave_gen_inst/_0687_ ),
    .B1_N(\wave_gen_inst/_1003_ ),
    .Y(\wave_gen_inst/_1004_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/_3881_  (.A1(\wave_gen_inst/_0987_ ),
    .A2(\wave_gen_inst/_0989_ ),
    .B1_N(\wave_gen_inst/_0985_ ),
    .Y(\wave_gen_inst/_1005_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3882_  (.A(\wave_gen_inst/counter[6] ),
    .B(net163),
    .Y(\wave_gen_inst/_1006_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3883_  (.A1(\wave_gen_inst/_1005_ ),
    .A2(\wave_gen_inst/_1006_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1007_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3884_  (.A1(\wave_gen_inst/_1005_ ),
    .A2(\wave_gen_inst/_1006_ ),
    .B1(\wave_gen_inst/_1007_ ),
    .Y(\wave_gen_inst/_1008_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3885_  (.A(net141),
    .B(\wave_gen_inst/_1002_ ),
    .C(\wave_gen_inst/_1004_ ),
    .D(\wave_gen_inst/_1008_ ),
    .Y(\wave_gen_inst/_1009_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/_3886_  (.A1(\wave_gen_inst/_0135_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_0997_ ),
    .B2(\wave_gen_inst/_1009_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0036_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3887_  (.A(\wave_gen_inst/_0685_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_1010_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3888_  (.A1(\wave_gen_inst/param1[7] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_1010_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_1011_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3889_  (.A1(\wave_gen_inst/sign ),
    .A2(\wave_gen_inst/_0780_ ),
    .A3(\wave_gen_inst/_0822_ ),
    .B1(\wave_gen_inst/_1011_ ),
    .Y(\wave_gen_inst/_1012_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3890_  (.A(\wave_gen_inst/_0133_ ),
    .B(\wave_gen_inst/_1000_ ),
    .Y(\wave_gen_inst/_1013_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3891_  (.A(net163),
    .B(\wave_gen_inst/_0685_ ),
    .Y(\wave_gen_inst/_1014_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3892_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0780_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1015_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3893_  (.A(\wave_gen_inst/_1014_ ),
    .B(\wave_gen_inst/_1015_ ),
    .Y(\wave_gen_inst/_1016_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3894_  (.A(\wave_gen_inst/counter[6] ),
    .B(net163),
    .Y(\wave_gen_inst/_1017_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3895_  (.A(\wave_gen_inst/counter[6] ),
    .B(net163),
    .Y(\wave_gen_inst/_1018_ ));
 sky130_fd_sc_hd__o311a_1 \wave_gen_inst/_3896_  (.A1(\wave_gen_inst/_0966_ ),
    .A2(\wave_gen_inst/_0986_ ),
    .A3(\wave_gen_inst/_0988_ ),
    .B1(\wave_gen_inst/_1018_ ),
    .C1(\wave_gen_inst/_0985_ ),
    .X(\wave_gen_inst/_1019_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3897_  (.A(\wave_gen_inst/counter[7] ),
    .B(net163),
    .X(\wave_gen_inst/_1020_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_3898_  (.A(\wave_gen_inst/_1020_ ),
    .Y(\wave_gen_inst/_1021_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3899_  (.A1(\wave_gen_inst/_1017_ ),
    .A2(\wave_gen_inst/_1019_ ),
    .B1(\wave_gen_inst/_1021_ ),
    .Y(\wave_gen_inst/_1022_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3900_  (.A(\wave_gen_inst/_1017_ ),
    .B(\wave_gen_inst/_1021_ ),
    .C(\wave_gen_inst/_1019_ ),
    .X(\wave_gen_inst/_1023_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3901_  (.A(\wave_gen_inst/_0106_ ),
    .B(\wave_gen_inst/_1022_ ),
    .C(\wave_gen_inst/_1023_ ),
    .Y(\wave_gen_inst/_1024_ ));
 sky130_fd_sc_hd__o2111ai_1 \wave_gen_inst/_3902_  (.A1(\wave_gen_inst/_0919_ ),
    .A2(\wave_gen_inst/_1013_ ),
    .B1(\wave_gen_inst/_1016_ ),
    .C1(\wave_gen_inst/_1024_ ),
    .D1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1025_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3903_  (.A1(\wave_gen_inst/_1753_ ),
    .A2(\wave_gen_inst/_1012_ ),
    .B1(\wave_gen_inst/_1025_ ),
    .Y(\wave_gen_inst/_1026_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3904_  (.A1(\wave_gen_inst/_0133_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_1026_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0037_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3905_  (.A(\wave_gen_inst/_0680_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_1027_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3906_  (.A1(\wave_gen_inst/param1[8] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_1027_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_1028_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_3907_  (.A1(\wave_gen_inst/sign ),
    .A2(\wave_gen_inst/_0777_ ),
    .A3(\wave_gen_inst/_0822_ ),
    .B1(\wave_gen_inst/_1028_ ),
    .Y(\wave_gen_inst/_1029_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3908_  (.A(\wave_gen_inst/_1753_ ),
    .B(\wave_gen_inst/_1029_ ),
    .Y(\wave_gen_inst/_1030_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3909_  (.A(net163),
    .B(\wave_gen_inst/_0680_ ),
    .Y(\wave_gen_inst/_1031_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3911_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0777_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1033_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3912_  (.A(\wave_gen_inst/_0133_ ),
    .B(\wave_gen_inst/_1000_ ),
    .Y(\wave_gen_inst/_1034_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3913_  (.A(\wave_gen_inst/counter[8] ),
    .B(\wave_gen_inst/_1034_ ),
    .Y(\wave_gen_inst/_1035_ ));
 sky130_fd_sc_hd__nor3_2 \wave_gen_inst/_3914_  (.A(\wave_gen_inst/_0133_ ),
    .B(\wave_gen_inst/_1590_ ),
    .C(\wave_gen_inst/_1000_ ),
    .Y(\wave_gen_inst/_1036_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3915_  (.A(\wave_gen_inst/_0919_ ),
    .B(\wave_gen_inst/_1035_ ),
    .C(\wave_gen_inst/_1036_ ),
    .Y(\wave_gen_inst/_1037_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3916_  (.A(\wave_gen_inst/counter[7] ),
    .B(net163),
    .Y(\wave_gen_inst/_1038_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3917_  (.A(\wave_gen_inst/_1038_ ),
    .B(\wave_gen_inst/_1023_ ),
    .Y(\wave_gen_inst/_1039_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3918_  (.A(\wave_gen_inst/counter[8] ),
    .B(net163),
    .X(\wave_gen_inst/_1040_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3919_  (.A(\wave_gen_inst/_1039_ ),
    .B(\wave_gen_inst/_1040_ ),
    .Y(\wave_gen_inst/_1041_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3920_  (.A1(\wave_gen_inst/_0111_ ),
    .A2(\wave_gen_inst/_1041_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1042_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3921_  (.A1(\wave_gen_inst/_1031_ ),
    .A2(\wave_gen_inst/_1033_ ),
    .B1(\wave_gen_inst/_1037_ ),
    .C1(\wave_gen_inst/_1042_ ),
    .Y(\wave_gen_inst/_1043_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/_3922_  (.A1(\wave_gen_inst/_1590_ ),
    .A2(net141),
    .B1(\wave_gen_inst/_1030_ ),
    .B2(\wave_gen_inst/_1043_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0038_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3923_  (.A(\wave_gen_inst/_0679_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_1044_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3924_  (.A1(\wave_gen_inst/param1[9] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_1044_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_1045_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3925_  (.A(\wave_gen_inst/sign ),
    .B(\wave_gen_inst/_0775_ ),
    .C(\wave_gen_inst/_0822_ ),
    .X(\wave_gen_inst/_1046_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3926_  (.A1(\wave_gen_inst/_1045_ ),
    .A2(\wave_gen_inst/_1046_ ),
    .B1(\wave_gen_inst/_0944_ ),
    .Y(\wave_gen_inst/_1047_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3927_  (.A(net163),
    .B(\wave_gen_inst/_0679_ ),
    .Y(\wave_gen_inst/_1048_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3928_  (.A(\wave_gen_inst/_0970_ ),
    .B(\wave_gen_inst/_1048_ ),
    .Y(\wave_gen_inst/_1049_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3929_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0775_ ),
    .B1(\wave_gen_inst/_1049_ ),
    .Y(\wave_gen_inst/_1050_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3930_  (.A(\wave_gen_inst/counter[9] ),
    .B(\wave_gen_inst/_1036_ ),
    .Y(\wave_gen_inst/_1051_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_3931_  (.A(net829),
    .B(\wave_gen_inst/_1036_ ),
    .Y(\wave_gen_inst/_1052_ ));
 sky130_fd_sc_hd__nor3b_1 \wave_gen_inst/_3932_  (.A(\wave_gen_inst/_0919_ ),
    .B(\wave_gen_inst/_1051_ ),
    .C_N(\wave_gen_inst/_1052_ ),
    .Y(\wave_gen_inst/_1053_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3933_  (.A(\wave_gen_inst/counter[9] ),
    .B(net163),
    .X(\wave_gen_inst/_1054_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3934_  (.A1(\wave_gen_inst/_1590_ ),
    .A2(\wave_gen_inst/_0232_ ),
    .B1(\wave_gen_inst/_1038_ ),
    .C1(\wave_gen_inst/_1023_ ),
    .Y(\wave_gen_inst/_1055_ ));
 sky130_fd_sc_hd__o211a_2 \wave_gen_inst/_3935_  (.A1(\wave_gen_inst/counter[8] ),
    .A2(net163),
    .B1(\wave_gen_inst/_1054_ ),
    .C1(\wave_gen_inst/_1055_ ),
    .X(\wave_gen_inst/_1056_ ));
 sky130_fd_sc_hd__a21boi_0 \wave_gen_inst/_3936_  (.A1(\wave_gen_inst/_1590_ ),
    .A2(\wave_gen_inst/_0232_ ),
    .B1_N(\wave_gen_inst/_1055_ ),
    .Y(\wave_gen_inst/_1057_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3937_  (.A1(\wave_gen_inst/_1054_ ),
    .A2(\wave_gen_inst/_1057_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1058_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3938_  (.A1(\wave_gen_inst/_1056_ ),
    .A2(\wave_gen_inst/_1058_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1059_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_3939_  (.A(\wave_gen_inst/_1047_ ),
    .B(\wave_gen_inst/_1050_ ),
    .C(\wave_gen_inst/_1053_ ),
    .D(\wave_gen_inst/_1059_ ),
    .Y(\wave_gen_inst/_1060_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3940_  (.A1(\wave_gen_inst/_1646_ ),
    .A2(\wave_gen_inst/_0602_ ),
    .B1(\wave_gen_inst/_1060_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0039_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3941_  (.A1(\wave_gen_inst/param1[10] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_1061_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3942_  (.A1(\wave_gen_inst/_0674_ ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_1061_ ),
    .Y(\wave_gen_inst/_1062_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3943_  (.A(\wave_gen_inst/sign ),
    .B(\wave_gen_inst/_0774_ ),
    .C(\wave_gen_inst/_0822_ ),
    .Y(\wave_gen_inst/_1063_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3944_  (.A1(\wave_gen_inst/_1062_ ),
    .A2(\wave_gen_inst/_1063_ ),
    .B1(\wave_gen_inst/_1753_ ),
    .Y(\wave_gen_inst/_1064_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3945_  (.A(net163),
    .B(\wave_gen_inst/_0674_ ),
    .Y(\wave_gen_inst/_1065_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3947_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0774_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1067_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3948_  (.A(\wave_gen_inst/_0123_ ),
    .B(\wave_gen_inst/_1052_ ),
    .Y(\wave_gen_inst/_1068_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3949_  (.A1(\wave_gen_inst/counter[9] ),
    .A2(net163),
    .B1(\wave_gen_inst/_1056_ ),
    .Y(\wave_gen_inst/_1069_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3950_  (.A(\wave_gen_inst/counter[10] ),
    .B(net163),
    .Y(\wave_gen_inst/_1070_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3951_  (.A1(\wave_gen_inst/_1069_ ),
    .A2(\wave_gen_inst/_1070_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1071_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3952_  (.A1(\wave_gen_inst/_1069_ ),
    .A2(\wave_gen_inst/_1070_ ),
    .B1(\wave_gen_inst/_1071_ ),
    .Y(\wave_gen_inst/_1072_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3953_  (.A(\wave_gen_inst/_0602_ ),
    .B(\wave_gen_inst/_1072_ ),
    .Y(\wave_gen_inst/_1073_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3954_  (.A1(\wave_gen_inst/_0919_ ),
    .A2(\wave_gen_inst/_1068_ ),
    .B1(\wave_gen_inst/_1073_ ),
    .Y(\wave_gen_inst/_1074_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3955_  (.A1(\wave_gen_inst/_1065_ ),
    .A2(\wave_gen_inst/_1067_ ),
    .B1(\wave_gen_inst/_1074_ ),
    .Y(\wave_gen_inst/_1075_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/_3956_  (.A1(\wave_gen_inst/_0123_ ),
    .A2(\wave_gen_inst/_0602_ ),
    .B1(\wave_gen_inst/_1064_ ),
    .B2(\wave_gen_inst/_1075_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0040_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3957_  (.A(\wave_gen_inst/_0232_ ),
    .B(\wave_gen_inst/_0773_ ),
    .Y(\wave_gen_inst/_1076_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3958_  (.A1(net163),
    .A2(\wave_gen_inst/_0672_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1077_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_3959_  (.A1(net829),
    .A2(\wave_gen_inst/counter[10] ),
    .A3(\wave_gen_inst/_1036_ ),
    .B1(\wave_gen_inst/counter[11] ),
    .Y(\wave_gen_inst/_1078_ ));
 sky130_fd_sc_hd__nor3_4 \wave_gen_inst/_3960_  (.A(\wave_gen_inst/_0123_ ),
    .B(\wave_gen_inst/_0124_ ),
    .C(\wave_gen_inst/_1052_ ),
    .Y(\wave_gen_inst/_1079_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3961_  (.A(\wave_gen_inst/counter[10] ),
    .B(net163),
    .X(\wave_gen_inst/_1080_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3962_  (.A(\wave_gen_inst/_1056_ ),
    .B(\wave_gen_inst/_1080_ ),
    .Y(\wave_gen_inst/_1081_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_3963_  (.A1(net959),
    .A2(net943),
    .B1(net163),
    .Y(\wave_gen_inst/_1082_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3964_  (.A(\wave_gen_inst/_1081_ ),
    .B(\wave_gen_inst/_1082_ ),
    .Y(\wave_gen_inst/_1083_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3965_  (.A(\wave_gen_inst/counter[11] ),
    .B(net163),
    .X(\wave_gen_inst/_1084_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3966_  (.A1(\wave_gen_inst/_1083_ ),
    .A2(\wave_gen_inst/_1084_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_1085_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3967_  (.A1(\wave_gen_inst/_1083_ ),
    .A2(\wave_gen_inst/_1084_ ),
    .B1(\wave_gen_inst/_1085_ ),
    .Y(\wave_gen_inst/_1086_ ));
 sky130_fd_sc_hd__o311ai_1 \wave_gen_inst/_3968_  (.A1(\wave_gen_inst/_0919_ ),
    .A2(net830),
    .A3(\wave_gen_inst/_1079_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .C1(\wave_gen_inst/_1086_ ),
    .Y(\wave_gen_inst/_1087_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3969_  (.A(\wave_gen_inst/_0672_ ),
    .B(\wave_gen_inst/_0718_ ),
    .Y(\wave_gen_inst/_1088_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3970_  (.A1(\wave_gen_inst/param1[11] ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_1088_ ),
    .C1(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_1089_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_3971_  (.A(\wave_gen_inst/sign ),
    .B(\wave_gen_inst/_0773_ ),
    .C(\wave_gen_inst/_0822_ ),
    .X(\wave_gen_inst/_1090_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3972_  (.A1(\wave_gen_inst/_1089_ ),
    .A2(\wave_gen_inst/_1090_ ),
    .B1(\wave_gen_inst/_0944_ ),
    .Y(\wave_gen_inst/_1091_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3973_  (.A1(\wave_gen_inst/_1076_ ),
    .A2(\wave_gen_inst/_1077_ ),
    .B1(net831),
    .C1(\wave_gen_inst/_1091_ ),
    .Y(\wave_gen_inst/_1092_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_3974_  (.A1(\wave_gen_inst/_0124_ ),
    .A2(\wave_gen_inst/_0602_ ),
    .B1(net832),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0041_ ));
 sky130_fd_sc_hd__mux2i_1 \wave_gen_inst/_3976_  (.A0(\wave_gen_inst/_0714_ ),
    .A1(\wave_gen_inst/_0772_ ),
    .S(\wave_gen_inst/_0232_ ),
    .Y(\wave_gen_inst/_1094_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_3977_  (.A(\wave_gen_inst/_1083_ ),
    .B(\wave_gen_inst/_1084_ ),
    .Y(\wave_gen_inst/_1095_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3978_  (.A1(\wave_gen_inst/_0124_ ),
    .A2(\wave_gen_inst/_0232_ ),
    .B1(\wave_gen_inst/_1095_ ),
    .Y(\wave_gen_inst/_1096_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3979_  (.A(\wave_gen_inst/counter[12] ),
    .B(net163),
    .X(\wave_gen_inst/_1097_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_3980_  (.A(\wave_gen_inst/_1096_ ),
    .B(\wave_gen_inst/_1097_ ),
    .Y(\wave_gen_inst/_1098_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_8 \wave_gen_inst/_3981_  (.A(net13),
    .SLEEP(\wave_gen_inst/_0162_ ),
    .X(\wave_gen_inst/_1099_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3983_  (.A1(\wave_gen_inst/counter[12] ),
    .A2(\wave_gen_inst/_1079_ ),
    .B1(\wave_gen_inst/_1099_ ),
    .Y(\wave_gen_inst/_1101_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_3984_  (.A1(\wave_gen_inst/counter[12] ),
    .A2(\wave_gen_inst/_1079_ ),
    .B1(\wave_gen_inst/_1101_ ),
    .Y(\wave_gen_inst/_1102_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_3985_  (.A1(\wave_gen_inst/_0111_ ),
    .A2(\wave_gen_inst/_1098_ ),
    .B1(\wave_gen_inst/_1102_ ),
    .C1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1103_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3986_  (.A1(\wave_gen_inst/_0970_ ),
    .A2(\wave_gen_inst/_1094_ ),
    .B1(net847),
    .Y(\wave_gen_inst/_1104_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3987_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1105_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3988_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1104_ ),
    .C(\wave_gen_inst/_1105_ ),
    .Y(\wave_gen_inst/_0042_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_3989_  (.A(\wave_gen_inst/_1056_ ),
    .B(\wave_gen_inst/_1080_ ),
    .C(\wave_gen_inst/_1084_ ),
    .D(\wave_gen_inst/_1097_ ),
    .Y(\wave_gen_inst/_1106_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_3990_  (.A1(\wave_gen_inst/counter[11] ),
    .A2(\wave_gen_inst/counter[12] ),
    .B1(net163),
    .Y(\wave_gen_inst/_1107_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_3991_  (.A(\wave_gen_inst/_1082_ ),
    .B(\wave_gen_inst/_1106_ ),
    .C(\wave_gen_inst/_1107_ ),
    .Y(\wave_gen_inst/_1108_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_3992_  (.A(\wave_gen_inst/counter[13] ),
    .B(net163),
    .X(\wave_gen_inst/_1109_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3993_  (.A(\wave_gen_inst/counter[13] ),
    .B(net163),
    .Y(\wave_gen_inst/_1110_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_3994_  (.A(\wave_gen_inst/_1109_ ),
    .B(\wave_gen_inst/_1110_ ),
    .Y(\wave_gen_inst/_1111_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_3995_  (.A(\wave_gen_inst/_1108_ ),
    .B(\wave_gen_inst/_1111_ ),
    .X(\wave_gen_inst/_1112_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_3996_  (.A1(\wave_gen_inst/counter[12] ),
    .A2(\wave_gen_inst/_1079_ ),
    .B1(\wave_gen_inst/counter[13] ),
    .Y(\wave_gen_inst/_1113_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_3997_  (.A(\wave_gen_inst/counter[12] ),
    .B(\wave_gen_inst/counter[13] ),
    .C(\wave_gen_inst/_1079_ ),
    .X(\wave_gen_inst/_1114_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_3998_  (.A(\wave_gen_inst/_1099_ ),
    .B(\wave_gen_inst/_1113_ ),
    .C(\wave_gen_inst/_1114_ ),
    .Y(\wave_gen_inst/_1115_ ));
 sky130_fd_sc_hd__or2_1 \wave_gen_inst/_3999_  (.A(\wave_gen_inst/counter[13] ),
    .B(\wave_gen_inst/_0638_ ),
    .X(\wave_gen_inst/_1116_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4000_  (.A1(\wave_gen_inst/counter[13] ),
    .A2(\wave_gen_inst/_0638_ ),
    .B1(\wave_gen_inst/_0232_ ),
    .Y(\wave_gen_inst/_1117_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/_4001_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0771_ ),
    .B1(\wave_gen_inst/_1116_ ),
    .B2(\wave_gen_inst/_1117_ ),
    .C1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1118_ ));
 sky130_fd_sc_hd__a2111oi_0 \wave_gen_inst/_4002_  (.A1(\wave_gen_inst/_0106_ ),
    .A2(\wave_gen_inst/_1112_ ),
    .B1(\wave_gen_inst/_1115_ ),
    .C1(net140),
    .D1(\wave_gen_inst/_1118_ ),
    .Y(\wave_gen_inst/_1119_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4003_  (.A(\wave_gen_inst/counter[13] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1120_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4004_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1119_ ),
    .C(\wave_gen_inst/_1120_ ),
    .Y(\wave_gen_inst/_0043_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4006_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1116_ ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1122_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4007_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1116_ ),
    .B1(\wave_gen_inst/_1122_ ),
    .Y(\wave_gen_inst/_1123_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4008_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0770_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .C1(\wave_gen_inst/_1123_ ),
    .Y(\wave_gen_inst/_1124_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4009_  (.A1(\wave_gen_inst/_1108_ ),
    .A2(\wave_gen_inst/_1111_ ),
    .B1(\wave_gen_inst/_1109_ ),
    .Y(\wave_gen_inst/_1125_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4010_  (.A(\wave_gen_inst/counter[14] ),
    .B(net163),
    .Y(\wave_gen_inst/_1126_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4011_  (.A1(\wave_gen_inst/_1125_ ),
    .A2(\wave_gen_inst/_1126_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1127_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4012_  (.A1(\wave_gen_inst/_1125_ ),
    .A2(\wave_gen_inst/_1126_ ),
    .B1(\wave_gen_inst/_1127_ ),
    .Y(\wave_gen_inst/_1128_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4013_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1114_ ),
    .B1(\wave_gen_inst/_0166_ ),
    .Y(\wave_gen_inst/_1129_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4014_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1114_ ),
    .B1(\wave_gen_inst/_1129_ ),
    .Y(\wave_gen_inst/_1130_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4015_  (.A(net140),
    .B(\wave_gen_inst/_1124_ ),
    .C(\wave_gen_inst/_1128_ ),
    .D(\wave_gen_inst/_1130_ ),
    .Y(\wave_gen_inst/_1131_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4016_  (.A(\wave_gen_inst/counter[14] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1132_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4017_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1131_ ),
    .C(\wave_gen_inst/_1132_ ),
    .Y(\wave_gen_inst/_0044_ ));
 sky130_fd_sc_hd__a311o_1 \wave_gen_inst/_4018_  (.A1(\wave_gen_inst/_1082_ ),
    .A2(\wave_gen_inst/_1106_ ),
    .A3(\wave_gen_inst/_1107_ ),
    .B1(\wave_gen_inst/_1109_ ),
    .C1(\wave_gen_inst/_1110_ ),
    .X(\wave_gen_inst/_1133_ ));
 sky130_fd_sc_hd__or2_2 \wave_gen_inst/_4019_  (.A(\wave_gen_inst/_1133_ ),
    .B(\wave_gen_inst/_1126_ ),
    .X(\wave_gen_inst/_1134_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4020_  (.A1(\wave_gen_inst/counter[13] ),
    .A2(\wave_gen_inst/counter[14] ),
    .B1(net162),
    .Y(\wave_gen_inst/_1135_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_4021_  (.A(\wave_gen_inst/counter[15] ),
    .B(net162),
    .Y(\wave_gen_inst/_1136_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4022_  (.A1(\wave_gen_inst/_1134_ ),
    .A2(\wave_gen_inst/_1135_ ),
    .B1(\wave_gen_inst/_1136_ ),
    .Y(\wave_gen_inst/_1137_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_4023_  (.A(\wave_gen_inst/_1134_ ),
    .B(\wave_gen_inst/_1135_ ),
    .C(\wave_gen_inst/_1136_ ),
    .X(\wave_gen_inst/_1138_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4024_  (.A1(\wave_gen_inst/_0737_ ),
    .A2(\wave_gen_inst/_1079_ ),
    .B1(\wave_gen_inst/counter[15] ),
    .X(\wave_gen_inst/_1139_ ));
 sky130_fd_sc_hd__nand3_2 \wave_gen_inst/_4025_  (.A(\wave_gen_inst/counter[15] ),
    .B(\wave_gen_inst/_0737_ ),
    .C(\wave_gen_inst/_1079_ ),
    .Y(\wave_gen_inst/_1140_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4026_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1116_ ),
    .B1(\wave_gen_inst/counter[15] ),
    .Y(\wave_gen_inst/_1141_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4027_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0769_ ),
    .B1(\wave_gen_inst/_0970_ ),
    .Y(\wave_gen_inst/_1142_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4028_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0639_ ),
    .A3(\wave_gen_inst/_1141_ ),
    .B1(\wave_gen_inst/_1142_ ),
    .Y(\wave_gen_inst/_1143_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_4029_  (.A1(\wave_gen_inst/_0166_ ),
    .A2(\wave_gen_inst/_1139_ ),
    .A3(\wave_gen_inst/_1140_ ),
    .B1(net140),
    .C1(\wave_gen_inst/_1143_ ),
    .Y(\wave_gen_inst/_1144_ ));
 sky130_fd_sc_hd__o31a_1 \wave_gen_inst/_4030_  (.A1(\wave_gen_inst/_0111_ ),
    .A2(\wave_gen_inst/_1137_ ),
    .A3(\wave_gen_inst/_1138_ ),
    .B1(\wave_gen_inst/_1144_ ),
    .X(\wave_gen_inst/_1145_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4031_  (.A(\wave_gen_inst/counter[15] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1146_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4032_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1145_ ),
    .C(\wave_gen_inst/_1146_ ),
    .Y(\wave_gen_inst/_0045_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4033_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0765_ ),
    .B1(\wave_gen_inst/_0970_ ),
    .Y(\wave_gen_inst/_1147_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4034_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0654_ ),
    .B1(\wave_gen_inst/_1147_ ),
    .Y(\wave_gen_inst/_1148_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4035_  (.A1(\wave_gen_inst/counter[15] ),
    .A2(\wave_gen_inst/pp ),
    .B1(\wave_gen_inst/_1137_ ),
    .Y(\wave_gen_inst/_1149_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_4036_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1150_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4037_  (.A(\wave_gen_inst/_1149_ ),
    .B(\wave_gen_inst/_1150_ ),
    .Y(\wave_gen_inst/_1151_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4038_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_1140_ ),
    .X(\wave_gen_inst/_1152_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_4039_  (.A1(\wave_gen_inst/_0111_ ),
    .A2(\wave_gen_inst/_1151_ ),
    .B1(\wave_gen_inst/_1152_ ),
    .B2(\wave_gen_inst/_1099_ ),
    .Y(\wave_gen_inst/_1153_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4040_  (.A(net140),
    .B(\wave_gen_inst/_1148_ ),
    .C(\wave_gen_inst/_1153_ ),
    .Y(\wave_gen_inst/_1154_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4041_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1155_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4042_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1154_ ),
    .C(\wave_gen_inst/_1155_ ),
    .Y(\wave_gen_inst/_0046_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4043_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/counter[17] ),
    .C(\wave_gen_inst/_0639_ ),
    .Y(\wave_gen_inst/_1156_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_4044_  (.A1(\wave_gen_inst/counter[16] ),
    .A2(\wave_gen_inst/_0639_ ),
    .B1(\wave_gen_inst/counter[17] ),
    .X(\wave_gen_inst/_1157_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4045_  (.A1(\wave_gen_inst/_1156_ ),
    .A2(\wave_gen_inst/_1157_ ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1158_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4046_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0811_ ),
    .B1(\wave_gen_inst/_1158_ ),
    .Y(\wave_gen_inst/_1159_ ));
 sky130_fd_sc_hd__o41ai_2 \wave_gen_inst/_4047_  (.A1(\wave_gen_inst/counter[13] ),
    .A2(\wave_gen_inst/counter[14] ),
    .A3(\wave_gen_inst/counter[15] ),
    .A4(\wave_gen_inst/counter[16] ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1160_ ));
 sky130_fd_sc_hd__o31ai_4 \wave_gen_inst/_4048_  (.A1(\wave_gen_inst/_1134_ ),
    .A2(\wave_gen_inst/_1136_ ),
    .A3(\wave_gen_inst/_1150_ ),
    .B1(\wave_gen_inst/_1160_ ),
    .Y(\wave_gen_inst/_1161_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4049_  (.A(\wave_gen_inst/counter[17] ),
    .B(\wave_gen_inst/pp ),
    .X(\wave_gen_inst/_1162_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_4050_  (.A(\wave_gen_inst/_1161_ ),
    .B(\wave_gen_inst/_1162_ ),
    .X(\wave_gen_inst/_1163_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4051_  (.A1(\wave_gen_inst/_1161_ ),
    .A2(\wave_gen_inst/_1162_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1164_ ));
 sky130_fd_sc_hd__nand3_2 \wave_gen_inst/_4052_  (.A(\wave_gen_inst/counter[14] ),
    .B(\wave_gen_inst/counter[15] ),
    .C(\wave_gen_inst/_1114_ ),
    .Y(\wave_gen_inst/_1165_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/_4053_  (.A(\wave_gen_inst/counter[16] ),
    .SLEEP(\wave_gen_inst/_1165_ ),
    .X(\wave_gen_inst/_1166_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4054_  (.A1(\wave_gen_inst/counter[17] ),
    .A2(\wave_gen_inst/_1166_ ),
    .B1(\wave_gen_inst/_1099_ ),
    .Y(\wave_gen_inst/_1167_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4055_  (.A1(\wave_gen_inst/counter[17] ),
    .A2(\wave_gen_inst/_1166_ ),
    .B1(\wave_gen_inst/_1167_ ),
    .Y(\wave_gen_inst/_1168_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/_4056_  (.A1(\wave_gen_inst/_1163_ ),
    .A2(\wave_gen_inst/_1164_ ),
    .B1(\wave_gen_inst/_1168_ ),
    .C1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1169_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4057_  (.A1(\wave_gen_inst/_0970_ ),
    .A2(\wave_gen_inst/_1159_ ),
    .B1(\wave_gen_inst/_1169_ ),
    .Y(\wave_gen_inst/_1170_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4058_  (.A(\wave_gen_inst/counter[17] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1171_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4059_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1170_ ),
    .C(\wave_gen_inst/_1171_ ),
    .Y(\wave_gen_inst/_0047_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4061_  (.A(\wave_gen_inst/counter[18] ),
    .B(\wave_gen_inst/_1156_ ),
    .Y(\wave_gen_inst/_1173_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4062_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_1173_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1174_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4063_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0817_ ),
    .B1(\wave_gen_inst/_1174_ ),
    .Y(\wave_gen_inst/_1175_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4064_  (.A1(\wave_gen_inst/counter[17] ),
    .A2(\wave_gen_inst/pp ),
    .B1(\wave_gen_inst/_1163_ ),
    .Y(\wave_gen_inst/_1176_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4065_  (.A(\wave_gen_inst/counter[18] ),
    .B(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1177_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_4066_  (.A(\wave_gen_inst/_1177_ ),
    .Y(\wave_gen_inst/_1178_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4067_  (.A(\wave_gen_inst/_1176_ ),
    .B(\wave_gen_inst/_1178_ ),
    .Y(\wave_gen_inst/_1179_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4068_  (.A1(\wave_gen_inst/counter[17] ),
    .A2(\wave_gen_inst/_1166_ ),
    .B1(\wave_gen_inst/counter[18] ),
    .Y(\wave_gen_inst/_1180_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_4069_  (.A(\wave_gen_inst/_0760_ ),
    .B_N(\wave_gen_inst/_1166_ ),
    .Y(\wave_gen_inst/_1181_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4070_  (.A(\wave_gen_inst/_1099_ ),
    .B(\wave_gen_inst/_1180_ ),
    .C(\wave_gen_inst/_1181_ ),
    .Y(\wave_gen_inst/_1182_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4071_  (.A1(\wave_gen_inst/_0106_ ),
    .A2(\wave_gen_inst/_1179_ ),
    .B1(\wave_gen_inst/_1182_ ),
    .Y(\wave_gen_inst/_1183_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4072_  (.A(\wave_gen_inst/counter[18] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1184_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_4073_  (.A1(\wave_gen_inst/_0833_ ),
    .A2(\wave_gen_inst/_1175_ ),
    .A3(\wave_gen_inst/_1183_ ),
    .B1(\wave_gen_inst/_1184_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0048_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4074_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0764_ ),
    .B1(\wave_gen_inst/_0970_ ),
    .Y(\wave_gen_inst/_1185_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4075_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0650_ ),
    .B1(\wave_gen_inst/_1185_ ),
    .Y(\wave_gen_inst/_1186_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4076_  (.A(\wave_gen_inst/_1163_ ),
    .B(\wave_gen_inst/_1178_ ),
    .Y(\wave_gen_inst/_1187_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4077_  (.A(\wave_gen_inst/pp ),
    .B(\wave_gen_inst/_0154_ ),
    .Y(\wave_gen_inst/_1188_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4078_  (.A(\wave_gen_inst/_1187_ ),
    .B(\wave_gen_inst/_1188_ ),
    .Y(\wave_gen_inst/_1189_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4079_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/pp ),
    .X(\wave_gen_inst/_1190_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4080_  (.A1(\wave_gen_inst/_1189_ ),
    .A2(\wave_gen_inst/_1190_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1191_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4081_  (.A1(\wave_gen_inst/_1189_ ),
    .A2(\wave_gen_inst/_1190_ ),
    .B1(\wave_gen_inst/_1191_ ),
    .Y(\wave_gen_inst/_1192_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4082_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_1181_ ),
    .Y(\wave_gen_inst/_1193_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4083_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/counter[19] ),
    .Y(\wave_gen_inst/_1194_ ));
 sky130_fd_sc_hd__nor4b_4 \wave_gen_inst/_4084_  (.A(\wave_gen_inst/_0738_ ),
    .B(\wave_gen_inst/_0760_ ),
    .C(\wave_gen_inst/_1194_ ),
    .D_N(\wave_gen_inst/_1079_ ),
    .Y(\wave_gen_inst/_1195_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4085_  (.A(\wave_gen_inst/_1099_ ),
    .B(\wave_gen_inst/_1193_ ),
    .C(\wave_gen_inst/_1195_ ),
    .Y(\wave_gen_inst/_1196_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4086_  (.A(net140),
    .B(\wave_gen_inst/_1186_ ),
    .C(\wave_gen_inst/_1192_ ),
    .D(\wave_gen_inst/_1196_ ),
    .Y(\wave_gen_inst/_1197_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4087_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1198_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4088_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1197_ ),
    .C(\wave_gen_inst/_1198_ ),
    .Y(\wave_gen_inst/_0049_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_4089_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/pp ),
    .C(\wave_gen_inst/_1189_ ),
    .X(\wave_gen_inst/_1199_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4090_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/pp ),
    .X(\wave_gen_inst/_1200_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4091_  (.A1(\wave_gen_inst/_1199_ ),
    .A2(\wave_gen_inst/_1200_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_1201_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4092_  (.A1(\wave_gen_inst/_1199_ ),
    .A2(\wave_gen_inst/_1200_ ),
    .B1(\wave_gen_inst/_1201_ ),
    .Y(\wave_gen_inst/_1202_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4093_  (.A(\wave_gen_inst/_0232_ ),
    .B(\wave_gen_inst/_0810_ ),
    .Y(\wave_gen_inst/_1203_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4094_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0653_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1204_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4095_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/_1195_ ),
    .Y(\wave_gen_inst/_1205_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4096_  (.A1(\wave_gen_inst/_1099_ ),
    .A2(\wave_gen_inst/_1205_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1206_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4097_  (.A1(\wave_gen_inst/_1203_ ),
    .A2(\wave_gen_inst/_1204_ ),
    .B1(\wave_gen_inst/_1206_ ),
    .Y(\wave_gen_inst/_1207_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4098_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1208_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4099_  (.A1(\wave_gen_inst/_1202_ ),
    .A2(\wave_gen_inst/_1207_ ),
    .B1(\wave_gen_inst/_1208_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0050_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4100_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(\wave_gen_inst/_0645_ ),
    .B1(\wave_gen_inst/counter[21] ),
    .Y(\wave_gen_inst/_1209_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4101_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0646_ ),
    .A3(\wave_gen_inst/_1209_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1210_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4102_  (.A1(\wave_gen_inst/pp ),
    .A2(\wave_gen_inst/_0819_ ),
    .B1(\wave_gen_inst/_1210_ ),
    .Y(\wave_gen_inst/_1211_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4103_  (.A(\wave_gen_inst/_1190_ ),
    .B(\wave_gen_inst/_1200_ ),
    .Y(\wave_gen_inst/_1212_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_4104_  (.A1(\wave_gen_inst/counter[19] ),
    .A2(\wave_gen_inst/counter[20] ),
    .A3(\wave_gen_inst/_0154_ ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1213_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4105_  (.A1(\wave_gen_inst/_1187_ ),
    .A2(\wave_gen_inst/_1212_ ),
    .B1(\wave_gen_inst/_1213_ ),
    .Y(\wave_gen_inst/_1214_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4106_  (.A(\wave_gen_inst/counter[21] ),
    .B(\wave_gen_inst/pp ),
    .X(\wave_gen_inst/_1215_ ));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 \wave_gen_inst/_4107_  (.A(\wave_gen_inst/_1214_ ),
    .SLEEP_B(\wave_gen_inst/_1215_ ),
    .X(\wave_gen_inst/_1216_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4108_  (.A(\wave_gen_inst/_0111_ ),
    .B(\wave_gen_inst/_1216_ ),
    .Y(\wave_gen_inst/_1217_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4109_  (.A1(\wave_gen_inst/_1214_ ),
    .A2(\wave_gen_inst/_1215_ ),
    .B1(\wave_gen_inst/_1217_ ),
    .Y(\wave_gen_inst/_1218_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4110_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(\wave_gen_inst/_1195_ ),
    .B1(\wave_gen_inst/counter[21] ),
    .X(\wave_gen_inst/_1219_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4111_  (.A(\wave_gen_inst/counter[20] ),
    .B(\wave_gen_inst/counter[21] ),
    .C(\wave_gen_inst/_1195_ ),
    .Y(\wave_gen_inst/_1220_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4112_  (.A1(\wave_gen_inst/_0166_ ),
    .A2(\wave_gen_inst/_1219_ ),
    .A3(\wave_gen_inst/_1220_ ),
    .B1(net140),
    .Y(\wave_gen_inst/_1221_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4113_  (.A(\wave_gen_inst/counter[21] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1222_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_4114_  (.A1(\wave_gen_inst/_1211_ ),
    .A2(\wave_gen_inst/_1218_ ),
    .A3(\wave_gen_inst/_1221_ ),
    .B1(\wave_gen_inst/_1222_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0051_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4115_  (.A1(net162),
    .A2(\wave_gen_inst/_0648_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1223_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4116_  (.A1(net162),
    .A2(\wave_gen_inst/_0752_ ),
    .B1(\wave_gen_inst/_1223_ ),
    .Y(\wave_gen_inst/_1224_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4117_  (.A1(\wave_gen_inst/counter[21] ),
    .A2(\wave_gen_inst/pp ),
    .B1(\wave_gen_inst/_1216_ ),
    .X(\wave_gen_inst/_1225_ ));
 sky130_fd_sc_hd__xor2_2 \wave_gen_inst/_4118_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/pp ),
    .X(\wave_gen_inst/_1226_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4119_  (.A1(\wave_gen_inst/_1225_ ),
    .A2(\wave_gen_inst/_1226_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_1227_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4120_  (.A1(\wave_gen_inst/_1225_ ),
    .A2(\wave_gen_inst/_1226_ ),
    .B1(\wave_gen_inst/_1227_ ),
    .Y(\wave_gen_inst/_1228_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4121_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/_1220_ ),
    .Y(\wave_gen_inst/_1229_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4122_  (.A1(\wave_gen_inst/_0166_ ),
    .A2(\wave_gen_inst/_1229_ ),
    .B1(net140),
    .Y(\wave_gen_inst/_1230_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4123_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1231_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_4124_  (.A1(\wave_gen_inst/_1224_ ),
    .A2(\wave_gen_inst/_1228_ ),
    .A3(\wave_gen_inst/_1230_ ),
    .B1(\wave_gen_inst/_1231_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0052_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4125_  (.A(\wave_gen_inst/_1216_ ),
    .B(\wave_gen_inst/_1226_ ),
    .Y(\wave_gen_inst/_1232_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_4126_  (.A1(\wave_gen_inst/counter[21] ),
    .A2(\wave_gen_inst/counter[22] ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1233_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4127_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1234_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4128_  (.A1(\wave_gen_inst/_1232_ ),
    .A2(\wave_gen_inst/_1233_ ),
    .B1(\wave_gen_inst/_1234_ ),
    .X(\wave_gen_inst/_1235_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4129_  (.A1(\wave_gen_inst/_1232_ ),
    .A2(\wave_gen_inst/_1233_ ),
    .A3(\wave_gen_inst/_1234_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_1236_ ));
 sky130_fd_sc_hd__a41oi_1 \wave_gen_inst/_4130_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(\wave_gen_inst/counter[21] ),
    .A3(\wave_gen_inst/counter[22] ),
    .A4(\wave_gen_inst/_1195_ ),
    .B1(\wave_gen_inst/counter[23] ),
    .Y(\wave_gen_inst/_1237_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4131_  (.A(\wave_gen_inst/_0842_ ),
    .B(\wave_gen_inst/_1165_ ),
    .Y(\wave_gen_inst/_1238_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4132_  (.A1(net162),
    .A2(\wave_gen_inst/_0651_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1239_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4133_  (.A1(net162),
    .A2(\wave_gen_inst/_0806_ ),
    .B1(\wave_gen_inst/_1239_ ),
    .Y(\wave_gen_inst/_1240_ ));
 sky130_fd_sc_hd__o311ai_2 \wave_gen_inst/_4134_  (.A1(\wave_gen_inst/_1099_ ),
    .A2(\wave_gen_inst/_1237_ ),
    .A3(\wave_gen_inst/_1238_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .C1(\wave_gen_inst/_1240_ ),
    .Y(\wave_gen_inst/_1241_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4135_  (.A1(\wave_gen_inst/_1235_ ),
    .A2(\wave_gen_inst/_1236_ ),
    .B1(\wave_gen_inst/_1241_ ),
    .Y(\wave_gen_inst/_1242_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4136_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1243_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4137_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1242_ ),
    .C(\wave_gen_inst/_1243_ ),
    .Y(\wave_gen_inst/_0053_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4138_  (.A(net162),
    .B(\wave_gen_inst/_0655_ ),
    .Y(\wave_gen_inst/_1244_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4139_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0809_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1245_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_4140_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/_1238_ ),
    .X(\wave_gen_inst/_1246_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4141_  (.A1(\wave_gen_inst/counter[24] ),
    .A2(\wave_gen_inst/_1238_ ),
    .B1(\wave_gen_inst/_0166_ ),
    .Y(\wave_gen_inst/_1247_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4142_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1248_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4143_  (.A(\wave_gen_inst/_1248_ ),
    .B(\wave_gen_inst/_1235_ ),
    .Y(\wave_gen_inst/_1249_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4144_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/pp ),
    .X(\wave_gen_inst/_1250_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4145_  (.A1(\wave_gen_inst/_1249_ ),
    .A2(\wave_gen_inst/_1250_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1251_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4146_  (.A1(\wave_gen_inst/_1249_ ),
    .A2(\wave_gen_inst/_1250_ ),
    .B1(\wave_gen_inst/_1251_ ),
    .Y(\wave_gen_inst/_1252_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4147_  (.A(net140),
    .B(\wave_gen_inst/_1252_ ),
    .Y(\wave_gen_inst/_1253_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4148_  (.A1(\wave_gen_inst/_1246_ ),
    .A2(\wave_gen_inst/_1247_ ),
    .B1(\wave_gen_inst/_1253_ ),
    .Y(\wave_gen_inst/_1254_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4149_  (.A1(\wave_gen_inst/_1244_ ),
    .A2(\wave_gen_inst/_1245_ ),
    .B1(\wave_gen_inst/_1254_ ),
    .Y(\wave_gen_inst/_1255_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4150_  (.A(\wave_gen_inst/counter[24] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1256_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4151_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1255_ ),
    .C(\wave_gen_inst/_1256_ ),
    .Y(\wave_gen_inst/_0054_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4152_  (.A(\wave_gen_inst/_1216_ ),
    .B(\wave_gen_inst/_1226_ ),
    .C(\wave_gen_inst/_1250_ ),
    .Y(\wave_gen_inst/_1257_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4153_  (.A1(\wave_gen_inst/counter[23] ),
    .A2(\wave_gen_inst/counter[24] ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1258_ ));
 sky130_fd_sc_hd__o211ai_2 \wave_gen_inst/_4154_  (.A1(\wave_gen_inst/_1234_ ),
    .A2(\wave_gen_inst/_1257_ ),
    .B1(\wave_gen_inst/_1258_ ),
    .C1(\wave_gen_inst/_1233_ ),
    .Y(\wave_gen_inst/_1259_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4155_  (.A(\wave_gen_inst/counter[25] ),
    .B(net162),
    .X(\wave_gen_inst/_1260_ ));
 sky130_fd_sc_hd__and2_0 \wave_gen_inst/_4156_  (.A(\wave_gen_inst/_1259_ ),
    .B(\wave_gen_inst/_1260_ ),
    .X(\wave_gen_inst/_1261_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4157_  (.A1(\wave_gen_inst/_1259_ ),
    .A2(\wave_gen_inst/_1260_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1262_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4158_  (.A(\wave_gen_inst/_1261_ ),
    .B(\wave_gen_inst/_1262_ ),
    .Y(\wave_gen_inst/_1263_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4159_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/_0660_ ),
    .Y(\wave_gen_inst/_1264_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4160_  (.A(net162),
    .B(\wave_gen_inst/_0804_ ),
    .Y(\wave_gen_inst/_1265_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_4161_  (.A1(net162),
    .A2(\wave_gen_inst/_0642_ ),
    .A3(\wave_gen_inst/_1264_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .C1(\wave_gen_inst/_1265_ ),
    .Y(\wave_gen_inst/_1266_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4162_  (.A1(\wave_gen_inst/counter[25] ),
    .A2(\wave_gen_inst/_1246_ ),
    .B1(\wave_gen_inst/_0166_ ),
    .Y(\wave_gen_inst/_1267_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4163_  (.A1(\wave_gen_inst/counter[25] ),
    .A2(\wave_gen_inst/_1246_ ),
    .B1(\wave_gen_inst/_1267_ ),
    .Y(\wave_gen_inst/_1268_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4164_  (.A(net140),
    .B(\wave_gen_inst/_1263_ ),
    .C(\wave_gen_inst/_1266_ ),
    .D(\wave_gen_inst/_1268_ ),
    .Y(\wave_gen_inst/_1269_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4165_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1270_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4166_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1269_ ),
    .C(\wave_gen_inst/_1270_ ),
    .Y(\wave_gen_inst/_0055_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4167_  (.A1(\wave_gen_inst/counter[25] ),
    .A2(net162),
    .B1(\wave_gen_inst/_1261_ ),
    .Y(\wave_gen_inst/_1271_ ));
 sky130_fd_sc_hd__xnor2_2 \wave_gen_inst/_4168_  (.A(\wave_gen_inst/counter[26] ),
    .B(net162),
    .Y(\wave_gen_inst/_1272_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4169_  (.A1(\wave_gen_inst/_1271_ ),
    .A2(\wave_gen_inst/_1272_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1273_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4170_  (.A1(\wave_gen_inst/_1271_ ),
    .A2(\wave_gen_inst/_1272_ ),
    .B1(\wave_gen_inst/_1273_ ),
    .Y(\wave_gen_inst/_1274_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4171_  (.A(net162),
    .B(\wave_gen_inst/_0750_ ),
    .Y(\wave_gen_inst/_1275_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4172_  (.A1(\wave_gen_inst/counter[26] ),
    .A2(\wave_gen_inst/_0642_ ),
    .B1(net162),
    .Y(\wave_gen_inst/_1276_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4173_  (.A1(\wave_gen_inst/counter[26] ),
    .A2(\wave_gen_inst/_0642_ ),
    .B1(\wave_gen_inst/_1276_ ),
    .Y(\wave_gen_inst/_1277_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4174_  (.A(\wave_gen_inst/_0829_ ),
    .B(\wave_gen_inst/_1275_ ),
    .C(\wave_gen_inst/_1277_ ),
    .Y(\wave_gen_inst/_1278_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4175_  (.A1(net818),
    .A2(\wave_gen_inst/_1246_ ),
    .B1(\wave_gen_inst/counter[26] ),
    .Y(\wave_gen_inst/_1279_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_4176_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/counter[26] ),
    .C(\wave_gen_inst/_1246_ ),
    .X(\wave_gen_inst/_1280_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4177_  (.A(\wave_gen_inst/_1099_ ),
    .B(\wave_gen_inst/_1279_ ),
    .C(\wave_gen_inst/_1280_ ),
    .Y(\wave_gen_inst/_1281_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4178_  (.A(net140),
    .B(\wave_gen_inst/_1274_ ),
    .C(\wave_gen_inst/_1278_ ),
    .D(\wave_gen_inst/_1281_ ),
    .Y(\wave_gen_inst/_1282_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4179_  (.A(\wave_gen_inst/counter[26] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1283_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4180_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1282_ ),
    .C(\wave_gen_inst/_1283_ ),
    .Y(\wave_gen_inst/_0056_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4181_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0758_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1284_ ));
 sky130_fd_sc_hd__a21boi_0 \wave_gen_inst/_4182_  (.A1(net162),
    .A2(\wave_gen_inst/_0644_ ),
    .B1_N(\wave_gen_inst/_1284_ ),
    .Y(\wave_gen_inst/_1285_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_4183_  (.A1(\wave_gen_inst/counter[25] ),
    .A2(\wave_gen_inst/counter[26] ),
    .B1(net162),
    .X(\wave_gen_inst/_1286_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4184_  (.A(\wave_gen_inst/_1259_ ),
    .B(\wave_gen_inst/_1260_ ),
    .Y(\wave_gen_inst/_1287_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4185_  (.A(\wave_gen_inst/_1287_ ),
    .B(\wave_gen_inst/_1272_ ),
    .Y(\wave_gen_inst/_1288_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4186_  (.A(\wave_gen_inst/counter[27] ),
    .B(net162),
    .X(\wave_gen_inst/_1289_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4187_  (.A(\wave_gen_inst/_1286_ ),
    .B(\wave_gen_inst/_1288_ ),
    .C(\wave_gen_inst/_1289_ ),
    .Y(\wave_gen_inst/_1290_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4188_  (.A1(\wave_gen_inst/_1286_ ),
    .A2(\wave_gen_inst/_1288_ ),
    .B1(\wave_gen_inst/_1289_ ),
    .Y(\wave_gen_inst/_1291_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4189_  (.A(\wave_gen_inst/_0106_ ),
    .B(\wave_gen_inst/_1291_ ),
    .Y(\wave_gen_inst/_1292_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_4190_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_1280_ ),
    .X(\wave_gen_inst/_1293_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4191_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_1280_ ),
    .Y(\wave_gen_inst/_1294_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_4192_  (.A(\wave_gen_inst/_1099_ ),
    .B(\wave_gen_inst/_1293_ ),
    .C(\wave_gen_inst/_1294_ ),
    .X(\wave_gen_inst/_1295_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4193_  (.A1(\wave_gen_inst/_1290_ ),
    .A2(\wave_gen_inst/_1292_ ),
    .B1(\wave_gen_inst/_1295_ ),
    .Y(\wave_gen_inst/_1296_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4194_  (.A(net140),
    .B(\wave_gen_inst/_1285_ ),
    .C(\wave_gen_inst/_1296_ ),
    .Y(\wave_gen_inst/_1297_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4195_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1298_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4196_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1297_ ),
    .C(\wave_gen_inst/_1298_ ),
    .Y(\wave_gen_inst/_0057_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4197_  (.A(\wave_gen_inst/counter[27] ),
    .B(net162),
    .Y(\wave_gen_inst/_1299_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4198_  (.A(\wave_gen_inst/_1299_ ),
    .B(\wave_gen_inst/_1291_ ),
    .Y(\wave_gen_inst/_1300_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4199_  (.A(\wave_gen_inst/counter[28] ),
    .B(net162),
    .X(\wave_gen_inst/_1301_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4200_  (.A1(\wave_gen_inst/_1300_ ),
    .A2(\wave_gen_inst/_1301_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1302_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4201_  (.A1(\wave_gen_inst/_1300_ ),
    .A2(\wave_gen_inst/_1301_ ),
    .B1(\wave_gen_inst/_1302_ ),
    .Y(\wave_gen_inst/_1303_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4202_  (.A(net162),
    .B(\wave_gen_inst/_0815_ ),
    .Y(\wave_gen_inst/_1304_ ));
 sky130_fd_sc_hd__a311oi_2 \wave_gen_inst/_4203_  (.A1(net162),
    .A2(\wave_gen_inst/_0662_ ),
    .A3(\wave_gen_inst/_0663_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .C1(\wave_gen_inst/_1304_ ),
    .Y(\wave_gen_inst/_1305_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4204_  (.A1(\wave_gen_inst/counter[28] ),
    .A2(\wave_gen_inst/_1293_ ),
    .B1(\wave_gen_inst/_0166_ ),
    .Y(\wave_gen_inst/_1306_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4205_  (.A1(\wave_gen_inst/counter[28] ),
    .A2(\wave_gen_inst/_1293_ ),
    .B1(\wave_gen_inst/_1306_ ),
    .Y(\wave_gen_inst/_1307_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4206_  (.A(net140),
    .B(\wave_gen_inst/_1303_ ),
    .C(\wave_gen_inst/_1305_ ),
    .D(\wave_gen_inst/_1307_ ),
    .Y(\wave_gen_inst/_1308_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4207_  (.A(\wave_gen_inst/counter[28] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1309_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4208_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1308_ ),
    .C(\wave_gen_inst/_1309_ ),
    .Y(\wave_gen_inst/_0058_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4209_  (.A(\wave_gen_inst/_1289_ ),
    .B(\wave_gen_inst/_1301_ ),
    .Y(\wave_gen_inst/_1310_ ));
 sky130_fd_sc_hd__o41ai_1 \wave_gen_inst/_4210_  (.A1(\wave_gen_inst/counter[25] ),
    .A2(\wave_gen_inst/counter[26] ),
    .A3(\wave_gen_inst/counter[27] ),
    .A4(\wave_gen_inst/counter[28] ),
    .B1(net162),
    .Y(\wave_gen_inst/_1311_ ));
 sky130_fd_sc_hd__o31ai_2 \wave_gen_inst/_4211_  (.A1(\wave_gen_inst/_1287_ ),
    .A2(\wave_gen_inst/_1272_ ),
    .A3(\wave_gen_inst/_1310_ ),
    .B1(\wave_gen_inst/_1311_ ),
    .Y(\wave_gen_inst/_1312_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4212_  (.A(\wave_gen_inst/counter[29] ),
    .B(net162),
    .X(\wave_gen_inst/_1313_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4213_  (.A1(\wave_gen_inst/_1312_ ),
    .A2(\wave_gen_inst/_1313_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_1314_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4214_  (.A1(\wave_gen_inst/_1312_ ),
    .A2(\wave_gen_inst/_1313_ ),
    .B1(\wave_gen_inst/_1314_ ),
    .Y(\wave_gen_inst/_1315_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4215_  (.A1(\wave_gen_inst/counter[28] ),
    .A2(\wave_gen_inst/_1293_ ),
    .B1(\wave_gen_inst/counter[29] ),
    .Y(\wave_gen_inst/_1316_ ));
 sky130_fd_sc_hd__nor4_2 \wave_gen_inst/_4216_  (.A(\wave_gen_inst/_0842_ ),
    .B(\wave_gen_inst/_0843_ ),
    .C(\wave_gen_inst/_0753_ ),
    .D(\wave_gen_inst/_1140_ ),
    .Y(\wave_gen_inst/_1317_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4217_  (.A(\wave_gen_inst/counter[29] ),
    .B(\wave_gen_inst/_0662_ ),
    .Y(\wave_gen_inst/_1318_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4218_  (.A1(\wave_gen_inst/_0151_ ),
    .A2(\wave_gen_inst/_0159_ ),
    .A3(\wave_gen_inst/_0641_ ),
    .B1(\wave_gen_inst/_0232_ ),
    .Y(\wave_gen_inst/_1319_ ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/_4219_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0808_ ),
    .B1(\wave_gen_inst/_1318_ ),
    .B2(\wave_gen_inst/_1319_ ),
    .C1(\wave_gen_inst/_0829_ ),
    .X(\wave_gen_inst/_1320_ ));
 sky130_fd_sc_hd__o311a_1 \wave_gen_inst/_4220_  (.A1(\wave_gen_inst/_1099_ ),
    .A2(\wave_gen_inst/_1316_ ),
    .A3(\wave_gen_inst/_1317_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .C1(\wave_gen_inst/_1320_ ),
    .X(\wave_gen_inst/_1321_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4221_  (.A(\wave_gen_inst/counter[29] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1322_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4222_  (.A1(\wave_gen_inst/_1315_ ),
    .A2(\wave_gen_inst/_1321_ ),
    .B1(\wave_gen_inst/_1322_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0059_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4223_  (.A(\wave_gen_inst/counter[29] ),
    .B(\wave_gen_inst/counter[30] ),
    .C(\wave_gen_inst/_0662_ ),
    .Y(\wave_gen_inst/_1323_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4224_  (.A1(\wave_gen_inst/counter[29] ),
    .A2(\wave_gen_inst/_0662_ ),
    .B1(\wave_gen_inst/counter[30] ),
    .Y(\wave_gen_inst/_1324_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_4225_  (.A_N(\wave_gen_inst/_1323_ ),
    .B(\wave_gen_inst/_1324_ ),
    .C(net162),
    .Y(\wave_gen_inst/_1325_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4226_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0814_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1326_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4227_  (.A(\wave_gen_inst/counter[30] ),
    .B(\wave_gen_inst/_1317_ ),
    .Y(\wave_gen_inst/_1327_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4228_  (.A1(\wave_gen_inst/_1099_ ),
    .A2(\wave_gen_inst/_1327_ ),
    .B1(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1328_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_4229_  (.A(\wave_gen_inst/counter[29] ),
    .B(net162),
    .C(\wave_gen_inst/_1312_ ),
    .X(\wave_gen_inst/_1329_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4230_  (.A(\wave_gen_inst/counter[30] ),
    .B(net162),
    .X(\wave_gen_inst/_1330_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4231_  (.A1(\wave_gen_inst/_1329_ ),
    .A2(\wave_gen_inst/_1330_ ),
    .B1(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1331_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4232_  (.A1(\wave_gen_inst/_1329_ ),
    .A2(\wave_gen_inst/_1330_ ),
    .B1(\wave_gen_inst/_1331_ ),
    .Y(\wave_gen_inst/_1332_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4233_  (.A1(\wave_gen_inst/_1325_ ),
    .A2(\wave_gen_inst/_1326_ ),
    .B1(\wave_gen_inst/_1328_ ),
    .C1(\wave_gen_inst/_1332_ ),
    .Y(\wave_gen_inst/_1333_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4234_  (.A(\wave_gen_inst/counter[30] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1334_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4235_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1333_ ),
    .C(\wave_gen_inst/_1334_ ),
    .Y(\wave_gen_inst/_0060_ ));
 sky130_fd_sc_hd__mux2i_1 \wave_gen_inst/_4236_  (.A0(net162),
    .A1(\wave_gen_inst/counter[30] ),
    .S(\wave_gen_inst/_1329_ ),
    .Y(\wave_gen_inst/_1335_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4237_  (.A1(\wave_gen_inst/counter[30] ),
    .A2(net162),
    .B1(\wave_gen_inst/_1335_ ),
    .Y(\wave_gen_inst/_1336_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4238_  (.A1(\wave_gen_inst/counter[31] ),
    .A2(\wave_gen_inst/_1336_ ),
    .B1(\wave_gen_inst/_0111_ ),
    .Y(\wave_gen_inst/_1337_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4239_  (.A1(\wave_gen_inst/counter[31] ),
    .A2(\wave_gen_inst/_1336_ ),
    .B1(\wave_gen_inst/_1337_ ),
    .Y(\wave_gen_inst/_1338_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4240_  (.A(\wave_gen_inst/counter[31] ),
    .B(\wave_gen_inst/_1323_ ),
    .Y(\wave_gen_inst/_1339_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4241_  (.A1(net162),
    .A2(\wave_gen_inst/_1339_ ),
    .B1(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1340_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4242_  (.A1(net162),
    .A2(\wave_gen_inst/_0757_ ),
    .B1(\wave_gen_inst/_1340_ ),
    .Y(\wave_gen_inst/_1341_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4243_  (.A1(\wave_gen_inst/counter[30] ),
    .A2(\wave_gen_inst/_1317_ ),
    .B1(\wave_gen_inst/counter[31] ),
    .X(\wave_gen_inst/_1342_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_4244_  (.A_N(\wave_gen_inst/_0844_ ),
    .B(\wave_gen_inst/_1293_ ),
    .Y(\wave_gen_inst/_1343_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4245_  (.A1(\wave_gen_inst/_0166_ ),
    .A2(\wave_gen_inst/_1342_ ),
    .A3(\wave_gen_inst/_1343_ ),
    .B1(net140),
    .Y(\wave_gen_inst/_1344_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4246_  (.A(\wave_gen_inst/counter[31] ),
    .B(\wave_gen_inst/_0833_ ),
    .Y(\wave_gen_inst/_1345_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/_4247_  (.A1(\wave_gen_inst/_1338_ ),
    .A2(\wave_gen_inst/_1341_ ),
    .A3(\wave_gen_inst/_1344_ ),
    .B1(\wave_gen_inst/_1345_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0061_ ));
 sky130_fd_sc_hd__or3b_1 \wave_gen_inst/_4248_  (.A(\wave_gen_inst/param1[0] ),
    .B(\wave_gen_inst/_0718_ ),
    .C_N(\wave_gen_inst/sign ),
    .X(\wave_gen_inst/_1346_ ));
 sky130_fd_sc_hd__o21bai_1 \wave_gen_inst/_4249_  (.A1(\wave_gen_inst/_0699_ ),
    .A2(\wave_gen_inst/_0822_ ),
    .B1_N(\wave_gen_inst/sign ),
    .Y(\wave_gen_inst/_1347_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4250_  (.A1(\wave_gen_inst/_0699_ ),
    .A2(\wave_gen_inst/_0718_ ),
    .B1(\wave_gen_inst/_0944_ ),
    .Y(\wave_gen_inst/_1348_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4251_  (.A(\wave_gen_inst/_1346_ ),
    .B(\wave_gen_inst/_1347_ ),
    .C(\wave_gen_inst/_1348_ ),
    .Y(\wave_gen_inst/_1349_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4252_  (.A(\wave_gen_inst/counter[0] ),
    .B(\wave_gen_inst/_0919_ ),
    .Y(\wave_gen_inst/_1350_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4253_  (.A(\wave_gen_inst/_0699_ ),
    .B(\wave_gen_inst/_0829_ ),
    .Y(\wave_gen_inst/_1351_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4254_  (.A(\wave_gen_inst/_0106_ ),
    .B(net141),
    .C(\wave_gen_inst/_1350_ ),
    .D(\wave_gen_inst/_1351_ ),
    .Y(\wave_gen_inst/_1352_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4255_  (.A1(\wave_gen_inst/_0111_ ),
    .A2(\wave_gen_inst/_0833_ ),
    .B1(\wave_gen_inst/counter[0] ),
    .Y(\wave_gen_inst/_1353_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4256_  (.A1(\wave_gen_inst/_1349_ ),
    .A2(\wave_gen_inst/_1352_ ),
    .B1(\wave_gen_inst/_1353_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0063_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4257_  (.A(\wave_gen_inst/_2195_ ),
    .B(\wave_gen_inst/_0106_ ),
    .Y(\wave_gen_inst/_1354_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_4258_  (.A_N(net12),
    .B(net11),
    .Y(\wave_gen_inst/_1355_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_4259_  (.A(net13),
    .B(\wave_gen_inst/_0914_ ),
    .C(\wave_gen_inst/_1355_ ),
    .X(\wave_gen_inst/_1356_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4260_  (.A(net13),
    .B(\wave_gen_inst/_1762_ ),
    .Y(\wave_gen_inst/_1357_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4261_  (.A1(\wave_gen_inst/_1357_ ),
    .A2(\wave_gen_inst/_0164_ ),
    .B1(\wave_gen_inst/param1[0] ),
    .Y(\wave_gen_inst/_1358_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4262_  (.A(net13),
    .B(net15),
    .C(\wave_gen_inst/_1355_ ),
    .Y(\wave_gen_inst/_1359_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4263_  (.A1(\wave_gen_inst/counter[0] ),
    .A2(\wave_gen_inst/_0167_ ),
    .B1(\wave_gen_inst/_1359_ ),
    .Y(\wave_gen_inst/_1360_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_4264_  (.A(\wave_gen_inst/_1354_ ),
    .B(\wave_gen_inst/_1356_ ),
    .C(\wave_gen_inst/_1358_ ),
    .D(\wave_gen_inst/_1360_ ),
    .Y(\wave_gen_inst/_1361_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4265_  (.A(\wave_gen_inst/_0915_ ),
    .B(\wave_gen_inst/_1361_ ),
    .Y(\wave_gen_inst/_1362_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/_4266_  (.A(\wave_gen_inst/_0916_ ),
    .B_N(\wave_gen_inst/_1356_ ),
    .Y(\wave_gen_inst/_1363_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4267_  (.A(net15),
    .B(\wave_gen_inst/_1363_ ),
    .Y(\wave_gen_inst/_1364_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4268_  (.A(\wave_gen_inst/changed ),
    .B(\wave_gen_inst/_1362_ ),
    .C(\wave_gen_inst/_1364_ ),
    .Y(\wave_gen_inst/_0064_ ));
 sky130_fd_sc_hd__and4_1 \wave_gen_inst/_4269_  (.A(\wave_gen_inst/_1672_ ),
    .B(\wave_gen_inst/_0847_ ),
    .C(\wave_gen_inst/_0696_ ),
    .D(\wave_gen_inst/_0697_ ),
    .X(\wave_gen_inst/_1365_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_4270_  (.A(\wave_gen_inst/_0687_ ),
    .B(\wave_gen_inst/_0691_ ),
    .C(\wave_gen_inst/_0693_ ),
    .D(\wave_gen_inst/_1365_ ),
    .Y(\wave_gen_inst/_1366_ ));
 sky130_fd_sc_hd__and4b_1 \wave_gen_inst/_4271_  (.A_N(\wave_gen_inst/_1366_ ),
    .B(\wave_gen_inst/_0674_ ),
    .C(\wave_gen_inst/_0685_ ),
    .D(\wave_gen_inst/_0680_ ),
    .X(\wave_gen_inst/_1367_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/_4272_  (.A(\wave_gen_inst/_0679_ ),
    .B(\wave_gen_inst/_0672_ ),
    .C(\wave_gen_inst/_0715_ ),
    .D(\wave_gen_inst/_1367_ ),
    .Y(\wave_gen_inst/_1368_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_4273_  (.A1(\wave_gen_inst/_0659_ ),
    .A2(\wave_gen_inst/_0664_ ),
    .A3(\wave_gen_inst/_1368_ ),
    .B1(\wave_gen_inst/pp ),
    .Y(\wave_gen_inst/_1369_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \wave_gen_inst/_4274_  (.A1_N(\wave_gen_inst/_0232_ ),
    .A2_N(\wave_gen_inst/_0822_ ),
    .B1(\wave_gen_inst/_1369_ ),
    .B2(\wave_gen_inst/counter[31] ),
    .Y(\wave_gen_inst/_1370_ ));
 sky130_fd_sc_hd__nor4_2 \wave_gen_inst/_4275_  (.A(\wave_gen_inst/_1548_ ),
    .B(\wave_gen_inst/_1663_ ),
    .C(\wave_gen_inst/_1552_ ),
    .D(\wave_gen_inst/_1551_ ),
    .Y(\wave_gen_inst/_1371_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4276_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/param2[2] ),
    .C(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1372_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4277_  (.A(\wave_gen_inst/_1533_ ),
    .B(\wave_gen_inst/_0848_ ),
    .Y(\wave_gen_inst/_1373_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_4278_  (.A1(\wave_gen_inst/_1663_ ),
    .A2(\wave_gen_inst/_1705_ ),
    .B1(\wave_gen_inst/_1373_ ),
    .Y(\wave_gen_inst/_1374_ ));
 sky130_fd_sc_hd__a21boi_4 \wave_gen_inst/_4279_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1699_ ),
    .B1_N(\wave_gen_inst/_1374_ ),
    .Y(\wave_gen_inst/_1375_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/_4280_  (.A(\wave_gen_inst/_1372_ ),
    .B(\wave_gen_inst/_1375_ ),
    .X(\wave_gen_inst/_1376_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_4281_  (.A(\wave_gen_inst/_1526_ ),
    .B(\wave_gen_inst/_0848_ ),
    .Y(\wave_gen_inst/_1377_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4282_  (.A(\wave_gen_inst/_1721_ ),
    .B(\wave_gen_inst/_1377_ ),
    .Y(\wave_gen_inst/_1378_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4283_  (.A(\wave_gen_inst/_1372_ ),
    .B(\wave_gen_inst/_1375_ ),
    .Y(\wave_gen_inst/_1379_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_4284_  (.A(\wave_gen_inst/_1723_ ),
    .B(\wave_gen_inst/_1373_ ),
    .Y(\wave_gen_inst/_1380_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_4285_  (.A1(\wave_gen_inst/_1720_ ),
    .A2(\wave_gen_inst/_1377_ ),
    .B1(\wave_gen_inst/_1380_ ),
    .Y(\wave_gen_inst/_1381_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4286_  (.A1(\wave_gen_inst/_1601_ ),
    .A2(\wave_gen_inst/_1379_ ),
    .B1(\wave_gen_inst/_1381_ ),
    .X(\wave_gen_inst/_1382_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_4287_  (.A1(\wave_gen_inst/_1554_ ),
    .A2(\wave_gen_inst/_1371_ ),
    .B1(\wave_gen_inst/_1382_ ),
    .Y(\wave_gen_inst/_1383_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_4288_  (.A1(\wave_gen_inst/_1533_ ),
    .A2(\wave_gen_inst/_1572_ ),
    .B1(\wave_gen_inst/_1383_ ),
    .Y(\wave_gen_inst/_1384_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/_4289_  (.A(\wave_gen_inst/_1378_ ),
    .B(\wave_gen_inst/_1384_ ),
    .Y(\wave_gen_inst/_1385_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_4290_  (.A1(\wave_gen_inst/_1721_ ),
    .A2(\wave_gen_inst/_1376_ ),
    .B1(\wave_gen_inst/_1385_ ),
    .Y(\wave_gen_inst/_1386_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4291_  (.A1(\wave_gen_inst/counter[31] ),
    .A2(\wave_gen_inst/_1571_ ),
    .A3(\wave_gen_inst/_1371_ ),
    .B1(\wave_gen_inst/_1386_ ),
    .Y(\wave_gen_inst/_1387_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4292_  (.A1(\wave_gen_inst/_1721_ ),
    .A2(\wave_gen_inst/_1375_ ),
    .B1(\wave_gen_inst/_1385_ ),
    .Y(\wave_gen_inst/_1388_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4293_  (.A1(\wave_gen_inst/_1721_ ),
    .A2(\wave_gen_inst/_1374_ ),
    .B1(\wave_gen_inst/_1385_ ),
    .Y(\wave_gen_inst/_1389_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/_4294_  (.A1(\wave_gen_inst/counter[29] ),
    .A2(\wave_gen_inst/_1388_ ),
    .B1(\wave_gen_inst/_1389_ ),
    .B2(\wave_gen_inst/counter[28] ),
    .Y(\wave_gen_inst/_1390_ ));
 sky130_fd_sc_hd__o31ai_2 \wave_gen_inst/_4295_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1533_ ),
    .A3(\wave_gen_inst/_1572_ ),
    .B1(\wave_gen_inst/_1383_ ),
    .Y(\wave_gen_inst/_1391_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/_4296_  (.A1(\wave_gen_inst/_1572_ ),
    .A2(\wave_gen_inst/_1377_ ),
    .B1(\wave_gen_inst/_1383_ ),
    .Y(\wave_gen_inst/_1392_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4297_  (.A(\wave_gen_inst/param2[1] ),
    .B(\wave_gen_inst/_1541_ ),
    .Y(\wave_gen_inst/_1393_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/_4298_  (.A(\wave_gen_inst/_1663_ ),
    .B(\wave_gen_inst/_1699_ ),
    .Y(\wave_gen_inst/_1394_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/_4299_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1393_ ),
    .B1(\wave_gen_inst/_1394_ ),
    .Y(\wave_gen_inst/_1395_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/_4300_  (.A(\wave_gen_inst/_1395_ ),
    .Y(\wave_gen_inst/_1396_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4301_  (.A(\wave_gen_inst/_1572_ ),
    .B(\wave_gen_inst/_1396_ ),
    .Y(\wave_gen_inst/_1397_ ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/_4302_  (.A(\wave_gen_inst/counter[18] ),
    .B(\wave_gen_inst/_1392_ ),
    .C(\wave_gen_inst/_1397_ ),
    .X(\wave_gen_inst/_1398_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_4303_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_1391_ ),
    .C(\wave_gen_inst/_1398_ ),
    .X(\wave_gen_inst/_1399_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4304_  (.A(\wave_gen_inst/counter[19] ),
    .B(\wave_gen_inst/_1391_ ),
    .X(\wave_gen_inst/_1400_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4305_  (.A1(\wave_gen_inst/_1392_ ),
    .A2(\wave_gen_inst/_1397_ ),
    .B1(\wave_gen_inst/counter[18] ),
    .Y(\wave_gen_inst/_1401_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4306_  (.A(\wave_gen_inst/_1398_ ),
    .B(\wave_gen_inst/_1400_ ),
    .C(\wave_gen_inst/_1401_ ),
    .Y(\wave_gen_inst/_1402_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4307_  (.A(\wave_gen_inst/_1572_ ),
    .B(\wave_gen_inst/_1394_ ),
    .Y(\wave_gen_inst/_1403_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4308_  (.A1(\wave_gen_inst/_1392_ ),
    .A2(\wave_gen_inst/_1403_ ),
    .B1(\wave_gen_inst/counter[17] ),
    .Y(\wave_gen_inst/_1404_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_4309_  (.A1(\wave_gen_inst/counter[17] ),
    .A2(\wave_gen_inst/_1403_ ),
    .B1(\wave_gen_inst/counter[16] ),
    .X(\wave_gen_inst/_1405_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4310_  (.A(\wave_gen_inst/_1392_ ),
    .B(\wave_gen_inst/_1405_ ),
    .Y(\wave_gen_inst/_1406_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_4311_  (.A_N(\wave_gen_inst/_1402_ ),
    .B(\wave_gen_inst/_1404_ ),
    .C(\wave_gen_inst/_1406_ ),
    .Y(\wave_gen_inst/_1407_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/_4312_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_1384_ ),
    .X(\wave_gen_inst/_1408_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4313_  (.A(\wave_gen_inst/_1572_ ),
    .B(\wave_gen_inst/_1375_ ),
    .Y(\wave_gen_inst/_1409_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4314_  (.A1(\wave_gen_inst/_1392_ ),
    .A2(\wave_gen_inst/_1409_ ),
    .B1(\wave_gen_inst/counter[21] ),
    .Y(\wave_gen_inst/_1410_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4315_  (.A1(\wave_gen_inst/_1724_ ),
    .A2(\wave_gen_inst/_1379_ ),
    .B1(\wave_gen_inst/_1392_ ),
    .Y(\wave_gen_inst/_1411_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4316_  (.A(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/_1411_ ),
    .Y(\wave_gen_inst/_1412_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_4317_  (.A(\wave_gen_inst/_1408_ ),
    .B(\wave_gen_inst/_1410_ ),
    .C(\wave_gen_inst/_1412_ ),
    .X(\wave_gen_inst/_1413_ ));
 sky130_fd_sc_hd__o21bai_1 \wave_gen_inst/_4318_  (.A1(\wave_gen_inst/_1572_ ),
    .A2(\wave_gen_inst/_1374_ ),
    .B1_N(\wave_gen_inst/_1392_ ),
    .Y(\wave_gen_inst/_1414_ ));
 sky130_fd_sc_hd__o32ai_2 \wave_gen_inst/_4319_  (.A1(\wave_gen_inst/counter[21] ),
    .A2(\wave_gen_inst/_1392_ ),
    .A3(\wave_gen_inst/_1409_ ),
    .B1(\wave_gen_inst/_1414_ ),
    .B2(\wave_gen_inst/counter[20] ),
    .Y(\wave_gen_inst/_1415_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4320_  (.A1(\wave_gen_inst/counter[20] ),
    .A2(\wave_gen_inst/_1414_ ),
    .B1(\wave_gen_inst/_1415_ ),
    .Y(\wave_gen_inst/_1416_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4321_  (.A(\wave_gen_inst/_1413_ ),
    .B(\wave_gen_inst/_1416_ ),
    .Y(\wave_gen_inst/_1417_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4322_  (.A1(\wave_gen_inst/_1399_ ),
    .A2(\wave_gen_inst/_1407_ ),
    .B1(\wave_gen_inst/_1417_ ),
    .Y(\wave_gen_inst/_1418_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_4323_  (.A_N(\wave_gen_inst/counter[22] ),
    .B(\wave_gen_inst/_1411_ ),
    .Y(\wave_gen_inst/_1419_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_4324_  (.A(\wave_gen_inst/counter[23] ),
    .B(\wave_gen_inst/_1384_ ),
    .C(\wave_gen_inst/_1419_ ),
    .X(\wave_gen_inst/_1420_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4325_  (.A(\wave_gen_inst/counter[2] ),
    .B(\wave_gen_inst/_1723_ ),
    .C(\wave_gen_inst/_1395_ ),
    .Y(\wave_gen_inst/_1421_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4326_  (.A(\wave_gen_inst/param2[2] ),
    .B(\wave_gen_inst/_1533_ ),
    .C(\wave_gen_inst/_1705_ ),
    .Y(\wave_gen_inst/_1422_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4327_  (.A(\wave_gen_inst/_1723_ ),
    .B(\wave_gen_inst/_1422_ ),
    .Y(\wave_gen_inst/_1423_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4328_  (.A(\wave_gen_inst/_1655_ ),
    .B(\wave_gen_inst/_1423_ ),
    .Y(\wave_gen_inst/_1424_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4329_  (.A1(\wave_gen_inst/_1723_ ),
    .A2(\wave_gen_inst/_1395_ ),
    .B1(\wave_gen_inst/counter[2] ),
    .Y(\wave_gen_inst/_1425_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4330_  (.A(\wave_gen_inst/_1424_ ),
    .B(\wave_gen_inst/_1425_ ),
    .Y(\wave_gen_inst/_1426_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4331_  (.A(\wave_gen_inst/_1421_ ),
    .B(\wave_gen_inst/_1426_ ),
    .Y(\wave_gen_inst/_1427_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4332_  (.A(\wave_gen_inst/_1663_ ),
    .B(\wave_gen_inst/_1723_ ),
    .C(\wave_gen_inst/_1699_ ),
    .Y(\wave_gen_inst/_1428_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4333_  (.A(\wave_gen_inst/_1671_ ),
    .B(\wave_gen_inst/_1428_ ),
    .Y(\wave_gen_inst/_1429_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4334_  (.A1(\wave_gen_inst/counter[0] ),
    .A2(\wave_gen_inst/_0846_ ),
    .B1(\wave_gen_inst/_1427_ ),
    .C1(\wave_gen_inst/_1429_ ),
    .Y(\wave_gen_inst/_1430_ ));
 sky130_fd_sc_hd__nor3b_1 \wave_gen_inst/_4335_  (.A(\wave_gen_inst/counter[1] ),
    .B(\wave_gen_inst/_1427_ ),
    .C_N(\wave_gen_inst/_1428_ ),
    .Y(\wave_gen_inst/_1431_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_4336_  (.A(\wave_gen_inst/_1655_ ),
    .B(\wave_gen_inst/_1423_ ),
    .C(\wave_gen_inst/_1425_ ),
    .X(\wave_gen_inst/_1432_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4337_  (.A(\wave_gen_inst/_1555_ ),
    .B(\wave_gen_inst/_1375_ ),
    .Y(\wave_gen_inst/_1433_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4338_  (.A(\wave_gen_inst/counter[5] ),
    .B(\wave_gen_inst/_1433_ ),
    .Y(\wave_gen_inst/_1434_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4339_  (.A(\wave_gen_inst/_0135_ ),
    .B(\wave_gen_inst/_1555_ ),
    .C(\wave_gen_inst/_1376_ ),
    .Y(\wave_gen_inst/_1435_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4340_  (.A1(\wave_gen_inst/_1723_ ),
    .A2(\wave_gen_inst/_1379_ ),
    .B1(\wave_gen_inst/counter[6] ),
    .Y(\wave_gen_inst/_1436_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4341_  (.A(\wave_gen_inst/_0133_ ),
    .B(\wave_gen_inst/_1380_ ),
    .Y(\wave_gen_inst/_1437_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/_4342_  (.A(\wave_gen_inst/_1435_ ),
    .B(\wave_gen_inst/_1436_ ),
    .C(\wave_gen_inst/_1437_ ),
    .Y(\wave_gen_inst/_1438_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4343_  (.A(\wave_gen_inst/_1555_ ),
    .B(\wave_gen_inst/_1374_ ),
    .Y(\wave_gen_inst/_1439_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_4344_  (.A1(\wave_gen_inst/counter[5] ),
    .A2(\wave_gen_inst/_1433_ ),
    .B1(\wave_gen_inst/_1439_ ),
    .B2(\wave_gen_inst/counter[4] ),
    .Y(\wave_gen_inst/_1440_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4345_  (.A1(\wave_gen_inst/counter[4] ),
    .A2(\wave_gen_inst/_1439_ ),
    .B1(\wave_gen_inst/_1440_ ),
    .Y(\wave_gen_inst/_1441_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_4346_  (.A(\wave_gen_inst/_1434_ ),
    .B(\wave_gen_inst/_1438_ ),
    .C(\wave_gen_inst/_1441_ ),
    .X(\wave_gen_inst/_1442_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_4347_  (.A1(\wave_gen_inst/_1430_ ),
    .A2(\wave_gen_inst/_1431_ ),
    .A3(\wave_gen_inst/_1432_ ),
    .B1(\wave_gen_inst/_1442_ ),
    .Y(\wave_gen_inst/_1443_ ));
 sky130_fd_sc_hd__maj3_1 \wave_gen_inst/_4348_  (.A(\wave_gen_inst/_0133_ ),
    .B(\wave_gen_inst/_1380_ ),
    .C(\wave_gen_inst/_1436_ ),
    .X(\wave_gen_inst/_1444_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4349_  (.A1(\wave_gen_inst/_1434_ ),
    .A2(\wave_gen_inst/_1438_ ),
    .A3(\wave_gen_inst/_1440_ ),
    .B1(\wave_gen_inst/_1444_ ),
    .Y(\wave_gen_inst/_1445_ ));
 sky130_fd_sc_hd__o21bai_1 \wave_gen_inst/_4350_  (.A1(\wave_gen_inst/_1720_ ),
    .A2(\wave_gen_inst/_1375_ ),
    .B1_N(\wave_gen_inst/_1381_ ),
    .Y(\wave_gen_inst/_1446_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/_4351_  (.A1(\wave_gen_inst/_1554_ ),
    .A2(\wave_gen_inst/_1371_ ),
    .B1(\wave_gen_inst/_1382_ ),
    .X(\wave_gen_inst/_1447_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_4352_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1382_ ),
    .B1(\wave_gen_inst/_1447_ ),
    .B2(\wave_gen_inst/counter[15] ),
    .Y(\wave_gen_inst/_1448_ ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/_4353_  (.A1(\wave_gen_inst/counter[14] ),
    .A2(\wave_gen_inst/_1382_ ),
    .B1(\wave_gen_inst/_1447_ ),
    .B2(\wave_gen_inst/counter[15] ),
    .C1(\wave_gen_inst/_1448_ ),
    .X(\wave_gen_inst/_1449_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4354_  (.A1(\wave_gen_inst/counter[13] ),
    .A2(\wave_gen_inst/_1446_ ),
    .B1(\wave_gen_inst/_1449_ ),
    .Y(\wave_gen_inst/_1450_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4355_  (.A(\wave_gen_inst/_1720_ ),
    .B(\wave_gen_inst/_1374_ ),
    .Y(\wave_gen_inst/_1451_ ));
 sky130_fd_sc_hd__o32ai_2 \wave_gen_inst/_4356_  (.A1(\wave_gen_inst/counter[12] ),
    .A2(\wave_gen_inst/_1381_ ),
    .A3(\wave_gen_inst/_1451_ ),
    .B1(\wave_gen_inst/_1446_ ),
    .B2(\wave_gen_inst/counter[13] ),
    .Y(\wave_gen_inst/_1452_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/_4357_  (.A1(\wave_gen_inst/_1381_ ),
    .A2(\wave_gen_inst/_1451_ ),
    .B1(\wave_gen_inst/counter[12] ),
    .X(\wave_gen_inst/_1453_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4358_  (.A(\wave_gen_inst/_1452_ ),
    .B(\wave_gen_inst/_1453_ ),
    .Y(\wave_gen_inst/_1454_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4359_  (.A(\wave_gen_inst/_1450_ ),
    .B(\wave_gen_inst/_1454_ ),
    .Y(\wave_gen_inst/_1455_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4360_  (.A1(\wave_gen_inst/_1601_ ),
    .A2(\wave_gen_inst/_1395_ ),
    .B1(\wave_gen_inst/_1381_ ),
    .Y(\wave_gen_inst/_1456_ ));
 sky130_fd_sc_hd__xnor2_1 \wave_gen_inst/_4361_  (.A(\wave_gen_inst/_0123_ ),
    .B(\wave_gen_inst/_1456_ ),
    .Y(\wave_gen_inst/_1457_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/_4362_  (.A1(\wave_gen_inst/param2[2] ),
    .A2(\wave_gen_inst/_1533_ ),
    .A3(\wave_gen_inst/_1720_ ),
    .B1(\wave_gen_inst/_1380_ ),
    .Y(\wave_gen_inst/_1458_ ));
 sky130_fd_sc_hd__or2_0 \wave_gen_inst/_4363_  (.A(\wave_gen_inst/counter[11] ),
    .B(\wave_gen_inst/_1458_ ),
    .X(\wave_gen_inst/_1459_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4364_  (.A(\wave_gen_inst/counter[11] ),
    .B(\wave_gen_inst/_1458_ ),
    .Y(\wave_gen_inst/_1460_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4365_  (.A(\wave_gen_inst/_1720_ ),
    .B(\wave_gen_inst/_1394_ ),
    .Y(\wave_gen_inst/_1461_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4366_  (.A1(\wave_gen_inst/_1381_ ),
    .A2(\wave_gen_inst/_1461_ ),
    .B1(\wave_gen_inst/counter[9] ),
    .Y(\wave_gen_inst/_1462_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4367_  (.A(\wave_gen_inst/_1459_ ),
    .B(\wave_gen_inst/_1460_ ),
    .C(\wave_gen_inst/_1462_ ),
    .Y(\wave_gen_inst/_1463_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4368_  (.A(\wave_gen_inst/_1457_ ),
    .B(\wave_gen_inst/_1463_ ),
    .Y(\wave_gen_inst/_1464_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4369_  (.A1(\wave_gen_inst/counter[9] ),
    .A2(\wave_gen_inst/_1461_ ),
    .B1(\wave_gen_inst/counter[8] ),
    .Y(\wave_gen_inst/_1465_ ));
 sky130_fd_sc_hd__mux2i_1 \wave_gen_inst/_4370_  (.A0(\wave_gen_inst/_1465_ ),
    .A1(\wave_gen_inst/counter[8] ),
    .S(\wave_gen_inst/_1381_ ),
    .Y(\wave_gen_inst/_1466_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_4371_  (.A_N(\wave_gen_inst/_1455_ ),
    .B(\wave_gen_inst/_1464_ ),
    .C(\wave_gen_inst/_1466_ ),
    .Y(\wave_gen_inst/_1467_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4372_  (.A1(\wave_gen_inst/_1443_ ),
    .A2(\wave_gen_inst/_1445_ ),
    .B1(\wave_gen_inst/_1467_ ),
    .Y(\wave_gen_inst/_1468_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4373_  (.A(\wave_gen_inst/counter[15] ),
    .B(\wave_gen_inst/_1447_ ),
    .Y(\wave_gen_inst/_1469_ ));
 sky130_fd_sc_hd__nand3b_1 \wave_gen_inst/_4374_  (.A_N(\wave_gen_inst/_1381_ ),
    .B(\wave_gen_inst/_1464_ ),
    .C(\wave_gen_inst/_1465_ ),
    .Y(\wave_gen_inst/_1470_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4375_  (.A(\wave_gen_inst/_0123_ ),
    .B(\wave_gen_inst/_1456_ ),
    .C(\wave_gen_inst/_1460_ ),
    .Y(\wave_gen_inst/_1471_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/_4376_  (.A1(\wave_gen_inst/_1459_ ),
    .A2(\wave_gen_inst/_1470_ ),
    .A3(\wave_gen_inst/_1471_ ),
    .B1(\wave_gen_inst/_1455_ ),
    .Y(\wave_gen_inst/_1472_ ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/_4377_  (.A1(\wave_gen_inst/_1469_ ),
    .A2(\wave_gen_inst/_1448_ ),
    .B1(\wave_gen_inst/_1450_ ),
    .B2(\wave_gen_inst/_1452_ ),
    .C1(\wave_gen_inst/_1472_ ),
    .X(\wave_gen_inst/_1473_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4378_  (.A(\wave_gen_inst/counter[16] ),
    .B(\wave_gen_inst/_1392_ ),
    .Y(\wave_gen_inst/_1474_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4379_  (.A(\wave_gen_inst/_1474_ ),
    .B(\wave_gen_inst/_1404_ ),
    .Y(\wave_gen_inst/_1475_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4380_  (.A(\wave_gen_inst/_1406_ ),
    .B(\wave_gen_inst/_1402_ ),
    .C(\wave_gen_inst/_1417_ ),
    .D(\wave_gen_inst/_1475_ ),
    .Y(\wave_gen_inst/_1476_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4381_  (.A1(\wave_gen_inst/_1468_ ),
    .A2(\wave_gen_inst/_1473_ ),
    .B1(\wave_gen_inst/_1476_ ),
    .Y(\wave_gen_inst/_1477_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4382_  (.A(\wave_gen_inst/_1413_ ),
    .B(\wave_gen_inst/_1415_ ),
    .Y(\wave_gen_inst/_1478_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4383_  (.A(\wave_gen_inst/_1420_ ),
    .B(\wave_gen_inst/_1477_ ),
    .C(\wave_gen_inst/_1478_ ),
    .Y(\wave_gen_inst/_1479_ ));
 sky130_fd_sc_hd__or2_0 \wave_gen_inst/_4384_  (.A(\wave_gen_inst/_1378_ ),
    .B(\wave_gen_inst/_1384_ ),
    .X(\wave_gen_inst/_1480_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4385_  (.A1(\wave_gen_inst/_1721_ ),
    .A2(\wave_gen_inst/_1396_ ),
    .B1(\wave_gen_inst/_1385_ ),
    .Y(\wave_gen_inst/_1481_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4386_  (.A(\wave_gen_inst/param2[3] ),
    .B(\wave_gen_inst/_1571_ ),
    .C(\wave_gen_inst/_1422_ ),
    .Y(\wave_gen_inst/_1482_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4387_  (.A(\wave_gen_inst/_1385_ ),
    .B(\wave_gen_inst/_1482_ ),
    .Y(\wave_gen_inst/_1483_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_4388_  (.A1(\wave_gen_inst/counter[26] ),
    .A2(\wave_gen_inst/_1481_ ),
    .B1(\wave_gen_inst/_1483_ ),
    .B2(\wave_gen_inst/counter[27] ),
    .Y(\wave_gen_inst/_1484_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4389_  (.A(\wave_gen_inst/counter[26] ),
    .B(\wave_gen_inst/_1481_ ),
    .Y(\wave_gen_inst/_1485_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/_4390_  (.A1(\wave_gen_inst/_1721_ ),
    .A2(\wave_gen_inst/_1394_ ),
    .B1(\wave_gen_inst/_1385_ ),
    .Y(\wave_gen_inst/_1486_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4391_  (.A(\wave_gen_inst/counter[25] ),
    .B(\wave_gen_inst/_1486_ ),
    .Y(\wave_gen_inst/_1487_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/_4392_  (.A(\wave_gen_inst/counter[27] ),
    .B(\wave_gen_inst/_1483_ ),
    .Y(\wave_gen_inst/_1488_ ));
 sky130_fd_sc_hd__nand4b_1 \wave_gen_inst/_4393_  (.A_N(\wave_gen_inst/_1484_ ),
    .B(\wave_gen_inst/_1485_ ),
    .C(\wave_gen_inst/_1487_ ),
    .D(\wave_gen_inst/_1488_ ),
    .Y(\wave_gen_inst/_1489_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_4394_  (.A1(\wave_gen_inst/counter[24] ),
    .A2(\wave_gen_inst/_1480_ ),
    .B1(\wave_gen_inst/_1486_ ),
    .B2(\wave_gen_inst/counter[25] ),
    .Y(\wave_gen_inst/_1490_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4395_  (.A1(\wave_gen_inst/counter[24] ),
    .A2(\wave_gen_inst/_1480_ ),
    .B1(\wave_gen_inst/_1489_ ),
    .C1(\wave_gen_inst/_1490_ ),
    .Y(\wave_gen_inst/_1491_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4396_  (.A1(\wave_gen_inst/_1418_ ),
    .A2(\wave_gen_inst/_1479_ ),
    .B1(\wave_gen_inst/_1491_ ),
    .Y(\wave_gen_inst/_1492_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/_4397_  (.A_N(\wave_gen_inst/_1489_ ),
    .B(\wave_gen_inst/_1490_ ),
    .Y(\wave_gen_inst/_1493_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4398_  (.A(\wave_gen_inst/counter[28] ),
    .B(\wave_gen_inst/_1389_ ),
    .Y(\wave_gen_inst/_1494_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4399_  (.A1(\wave_gen_inst/_1484_ ),
    .A2(\wave_gen_inst/_1488_ ),
    .B1(\wave_gen_inst/_1494_ ),
    .Y(\wave_gen_inst/_1495_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/_4400_  (.A(\wave_gen_inst/_1492_ ),
    .B(\wave_gen_inst/_1493_ ),
    .C(\wave_gen_inst/_1495_ ),
    .Y(\wave_gen_inst/_1496_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/_4401_  (.A(\wave_gen_inst/counter[29] ),
    .B(\wave_gen_inst/_1388_ ),
    .Y(\wave_gen_inst/_1497_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/_4402_  (.A1(\wave_gen_inst/_1390_ ),
    .A2(\wave_gen_inst/_1496_ ),
    .B1(\wave_gen_inst/_1497_ ),
    .Y(\wave_gen_inst/_1498_ ));
 sky130_fd_sc_hd__o211ai_2 \wave_gen_inst/_4403_  (.A1(\wave_gen_inst/counter[0] ),
    .A2(\wave_gen_inst/_0846_ ),
    .B1(\wave_gen_inst/_1442_ ),
    .C1(\wave_gen_inst/_1430_ ),
    .Y(\wave_gen_inst/_1499_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4404_  (.A1(\wave_gen_inst/counter[29] ),
    .A2(\wave_gen_inst/_1388_ ),
    .B1(\wave_gen_inst/_1390_ ),
    .Y(\wave_gen_inst/_1500_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/_4405_  (.A(\wave_gen_inst/_1467_ ),
    .B(\wave_gen_inst/_1494_ ),
    .C(\wave_gen_inst/_1499_ ),
    .D(\wave_gen_inst/_1500_ ),
    .Y(\wave_gen_inst/_1501_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_4406_  (.A(\wave_gen_inst/_1491_ ),
    .B(\wave_gen_inst/_1476_ ),
    .C(\wave_gen_inst/_1501_ ),
    .X(\wave_gen_inst/_1502_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/_4407_  (.A1(\wave_gen_inst/counter[30] ),
    .A2(\wave_gen_inst/_1386_ ),
    .B1(\wave_gen_inst/_1498_ ),
    .B2(\wave_gen_inst/_1502_ ),
    .Y(\wave_gen_inst/_1503_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/_4408_  (.A1(\wave_gen_inst/_0152_ ),
    .A2(\wave_gen_inst/_1387_ ),
    .B1(\wave_gen_inst/_1503_ ),
    .Y(\wave_gen_inst/_1504_ ));
 sky130_fd_sc_hd__a211o_1 \wave_gen_inst/_4409_  (.A1(\wave_gen_inst/_1571_ ),
    .A2(\wave_gen_inst/_1371_ ),
    .B1(\wave_gen_inst/_1386_ ),
    .C1(\wave_gen_inst/counter[31] ),
    .X(\wave_gen_inst/_1505_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/_4410_  (.A(\wave_gen_inst/_0112_ ),
    .B(\wave_gen_inst/_1504_ ),
    .C(\wave_gen_inst/_1505_ ),
    .X(\wave_gen_inst/_1506_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/_4411_  (.A1(\wave_gen_inst/_0670_ ),
    .A2(net844),
    .B1(\wave_gen_inst/_0108_ ),
    .Y(\wave_gen_inst/_1507_ ));
 sky130_fd_sc_hd__a2111oi_0 \wave_gen_inst/_4412_  (.A1(\wave_gen_inst/_0111_ ),
    .A2(\wave_gen_inst/_1370_ ),
    .B1(\wave_gen_inst/_1506_ ),
    .C1(net845),
    .D1(\wave_gen_inst/_0969_ ),
    .Y(\wave_gen_inst/_1508_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/_4413_  (.A1(\wave_gen_inst/_0232_ ),
    .A2(\wave_gen_inst/_0969_ ),
    .B1(\wave_gen_inst/_1508_ ),
    .C1(\wave_gen_inst/changed ),
    .Y(\wave_gen_inst/_0065_ ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4414_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0000_ ),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4415_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0001_ ),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4416_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0002_ ),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4417_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0003_ ),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4418_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0004_ ),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4419_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0005_ ),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4420_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0006_ ),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4421_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0007_ ),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4422_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0008_ ),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4423_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0009_ ),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4424_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0010_ ),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4425_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0011_ ),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4426_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0012_ ),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4427_  (.CLK(clknet_leaf_74_clk),
    .D(\wave_gen_inst/_0013_ ),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4428_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0014_ ),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4429_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0015_ ),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4430_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0016_ ),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4431_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0017_ ),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4432_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0018_ ),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4433_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0019_ ),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4434_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0020_ ),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4435_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0021_ ),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4436_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0022_ ),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4437_  (.CLK(clknet_leaf_74_clk),
    .D(\wave_gen_inst/_0023_ ),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4438_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0024_ ),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4439_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0025_ ),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4440_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0026_ ),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4441_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0027_ ),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4442_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0028_ ),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4443_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0029_ ),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4444_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0030_ ),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4445_  (.CLK(clknet_leaf_66_clk),
    .D(\wave_gen_inst/_0031_ ),
    .Q(\wave_gen_inst/counter[1] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4446_  (.CLK(clknet_leaf_66_clk),
    .D(\wave_gen_inst/_0032_ ),
    .Q(\wave_gen_inst/counter[2] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4447_  (.CLK(clknet_leaf_66_clk),
    .D(\wave_gen_inst/_0033_ ),
    .Q(\wave_gen_inst/counter[3] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4448_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0034_ ),
    .Q(\wave_gen_inst/counter[4] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4449_  (.CLK(clknet_leaf_66_clk),
    .D(\wave_gen_inst/_0035_ ),
    .Q(\wave_gen_inst/counter[5] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4450_  (.CLK(clknet_leaf_66_clk),
    .D(\wave_gen_inst/_0036_ ),
    .Q(\wave_gen_inst/counter[6] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4451_  (.CLK(clknet_leaf_67_clk),
    .D(\wave_gen_inst/_0037_ ),
    .Q(\wave_gen_inst/counter[7] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4452_  (.CLK(clknet_leaf_67_clk),
    .D(\wave_gen_inst/_0038_ ),
    .Q(\wave_gen_inst/counter[8] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4453_  (.CLK(clknet_leaf_67_clk),
    .D(\wave_gen_inst/_0039_ ),
    .Q(\wave_gen_inst/counter[9] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4454_  (.CLK(clknet_leaf_67_clk),
    .D(\wave_gen_inst/_0040_ ),
    .Q(\wave_gen_inst/counter[10] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4455_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0041_ ),
    .Q(\wave_gen_inst/counter[11] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4456_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0042_ ),
    .Q(\wave_gen_inst/counter[12] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4457_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0043_ ),
    .Q(\wave_gen_inst/counter[13] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4458_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0044_ ),
    .Q(\wave_gen_inst/counter[14] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4459_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0045_ ),
    .Q(\wave_gen_inst/counter[15] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4460_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0046_ ),
    .Q(\wave_gen_inst/counter[16] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4461_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0047_ ),
    .Q(\wave_gen_inst/counter[17] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4462_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0048_ ),
    .Q(\wave_gen_inst/counter[18] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4463_  (.CLK(clknet_leaf_70_clk),
    .D(\wave_gen_inst/_0049_ ),
    .Q(\wave_gen_inst/counter[19] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4464_  (.CLK(clknet_leaf_70_clk),
    .D(\wave_gen_inst/_0050_ ),
    .Q(\wave_gen_inst/counter[20] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4465_  (.CLK(clknet_leaf_70_clk),
    .D(\wave_gen_inst/_0051_ ),
    .Q(\wave_gen_inst/counter[21] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4466_  (.CLK(clknet_leaf_70_clk),
    .D(\wave_gen_inst/_0052_ ),
    .Q(\wave_gen_inst/counter[22] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4467_  (.CLK(clknet_leaf_70_clk),
    .D(\wave_gen_inst/_0053_ ),
    .Q(\wave_gen_inst/counter[23] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4468_  (.CLK(clknet_leaf_69_clk),
    .D(\wave_gen_inst/_0054_ ),
    .Q(\wave_gen_inst/counter[24] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4469_  (.CLK(clknet_leaf_70_clk),
    .D(\wave_gen_inst/_0055_ ),
    .Q(\wave_gen_inst/counter[25] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4470_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0056_ ),
    .Q(\wave_gen_inst/counter[26] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4471_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0057_ ),
    .Q(\wave_gen_inst/counter[27] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4472_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0058_ ),
    .Q(\wave_gen_inst/counter[28] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4473_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0059_ ),
    .Q(\wave_gen_inst/counter[29] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4474_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0060_ ),
    .Q(\wave_gen_inst/counter[30] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4475_  (.CLK(clknet_leaf_73_clk),
    .D(\wave_gen_inst/_0061_ ),
    .Q(\wave_gen_inst/counter[31] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4476_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0062_ ),
    .Q(\wave_gen_inst/sign ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4477_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0063_ ),
    .Q(\wave_gen_inst/counter[0] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4478_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0064_ ),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4479_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0065_ ),
    .Q(\wave_gen_inst/pp ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4480_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0066_ ),
    .Q(\wave_gen_inst/param1[0] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4481_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0067_ ),
    .Q(\wave_gen_inst/param1[1] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4482_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0068_ ),
    .Q(\wave_gen_inst/param1[2] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4483_  (.CLK(clknet_leaf_65_clk),
    .D(\wave_gen_inst/_0069_ ),
    .Q(\wave_gen_inst/param1[3] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4484_  (.CLK(clknet_leaf_67_clk),
    .D(\wave_gen_inst/_0070_ ),
    .Q(\wave_gen_inst/param1[4] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4485_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0071_ ),
    .Q(\wave_gen_inst/param1[5] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4486_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0072_ ),
    .Q(\wave_gen_inst/param1[6] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4487_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0073_ ),
    .Q(\wave_gen_inst/param1[7] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4488_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0074_ ),
    .Q(\wave_gen_inst/param1[8] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4489_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0075_ ),
    .Q(\wave_gen_inst/param1[9] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4490_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0076_ ),
    .Q(\wave_gen_inst/param1[10] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4491_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0077_ ),
    .Q(\wave_gen_inst/param1[11] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4492_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0078_ ),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4493_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0079_ ),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4494_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0080_ ),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4495_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0081_ ),
    .Q(\wave_gen_inst/changed ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4496_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0082_ ),
    .Q(\wave_gen_inst/param1[0] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4497_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0083_ ),
    .Q(\wave_gen_inst/param1[1] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4498_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0084_ ),
    .Q(\wave_gen_inst/param1[2] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4499_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0085_ ),
    .Q(\wave_gen_inst/param1[3] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4500_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0086_ ),
    .Q(\wave_gen_inst/param1[4] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4501_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0087_ ),
    .Q(\wave_gen_inst/param1[5] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4502_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0088_ ),
    .Q(\wave_gen_inst/param1[6] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4503_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0089_ ),
    .Q(\wave_gen_inst/param1[7] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4504_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0090_ ),
    .Q(\wave_gen_inst/param1[8] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4505_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0091_ ),
    .Q(\wave_gen_inst/param1[9] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4506_  (.CLK(clknet_leaf_63_clk),
    .D(\wave_gen_inst/_0092_ ),
    .Q(\wave_gen_inst/param1[10] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4507_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0093_ ),
    .Q(\wave_gen_inst/param1[11] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4508_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0094_ ),
    .Q(\wave_gen_inst/param2[0] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4509_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0095_ ),
    .Q(\wave_gen_inst/param2[1] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4510_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0096_ ),
    .Q(\wave_gen_inst/param2[2] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4511_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0097_ ),
    .Q(\wave_gen_inst/param2[3] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4512_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0098_ ),
    .Q(\wave_gen_inst/param2[4] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4513_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0099_ ),
    .Q(\wave_gen_inst/param2[5] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4514_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0100_ ),
    .Q(\wave_gen_inst/param2[6] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4515_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0101_ ),
    .Q(\wave_gen_inst/param2[7] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4516_  (.CLK(clknet_leaf_62_clk),
    .D(\wave_gen_inst/_0102_ ),
    .Q(\wave_gen_inst/param2[8] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4517_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0103_ ),
    .Q(\wave_gen_inst/param2[9] ));
 sky130_fd_sc_hd__dfxtp_4 \wave_gen_inst/_4518_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0104_ ),
    .Q(\wave_gen_inst/param2[10] ));
 sky130_fd_sc_hd__dfxtp_2 \wave_gen_inst/_4519_  (.CLK(clknet_leaf_68_clk),
    .D(\wave_gen_inst/_0105_ ),
    .Q(\wave_gen_inst/param2[11] ));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_2738__473  (.HI(net473));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/rom/_247_  (.A_N(\wave_gen_inst/sine_phase[3] ),
    .B(\wave_gen_inst/sine_phase[0] ),
    .Y(\wave_gen_inst/rom/_166_ ));
 sky130_fd_sc_hd__xnor2_4 \wave_gen_inst/rom/_250_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_169_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \wave_gen_inst/rom/_252_  (.A1_N(\wave_gen_inst/sine_phase[1] ),
    .A2_N(\wave_gen_inst/rom/_166_ ),
    .B1(\wave_gen_inst/rom/_169_ ),
    .B2(\wave_gen_inst/sine_phase[3] ),
    .Y(\wave_gen_inst/rom/_171_ ));
 sky130_fd_sc_hd__nand2_4 \wave_gen_inst/rom/_256_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_175_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_259_  (.A1(\wave_gen_inst/sine_phase[1] ),
    .A2(\wave_gen_inst/rom/_175_ ),
    .B1(\wave_gen_inst/sine_phase[3] ),
    .Y(\wave_gen_inst/rom/_178_ ));
 sky130_fd_sc_hd__nand4b_1 \wave_gen_inst/rom/_260_  (.A_N(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/sine_phase[1] ),
    .D(\wave_gen_inst/sine_phase[3] ),
    .Y(\wave_gen_inst/rom/_179_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_261_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(\wave_gen_inst/rom/_179_ ),
    .Y(\wave_gen_inst/rom/_180_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/rom/_262_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_171_ ),
    .B1(\wave_gen_inst/rom/_178_ ),
    .B2(\wave_gen_inst/rom/_180_ ),
    .Y(\wave_gen_inst/rom/_181_ ));
 sky130_fd_sc_hd__lpflow_inputiso0n_1 \wave_gen_inst/rom/_263_  (.A(\wave_gen_inst/sine_phase[6] ),
    .SLEEP_B(\wave_gen_inst/rom/_181_ ),
    .X(\wave_gen_inst/rom/_182_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/rom/_265_  (.A(net70),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_184_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/rom/_266_  (.A(\wave_gen_inst/sine_phase[3] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_185_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_267_  (.A(\wave_gen_inst/rom/_169_ ),
    .B(\wave_gen_inst/rom/_185_ ),
    .Y(\wave_gen_inst/rom/_186_ ));
 sky130_fd_sc_hd__inv_6 \wave_gen_inst/rom/_268_  (.A(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_187_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_270_  (.A1(\wave_gen_inst/rom/_184_ ),
    .A2(\wave_gen_inst/rom/_186_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_189_ ));
 sky130_fd_sc_hd__inv_1 \wave_gen_inst/rom/_271_  (.A(\wave_gen_inst/sine_phase[0] ),
    .Y(\wave_gen_inst/rom/_190_ ));
 sky130_fd_sc_hd__nand2b_1 \wave_gen_inst/rom/_272_  (.A_N(\wave_gen_inst/sine_phase[1] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_191_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_273_  (.A(\wave_gen_inst/rom/_190_ ),
    .B(\wave_gen_inst/rom/_191_ ),
    .Y(\wave_gen_inst/rom/_192_ ));
 sky130_fd_sc_hd__nand2b_2 \wave_gen_inst/rom/_274_  (.A_N(\wave_gen_inst/sine_phase[4] ),
    .B(net70),
    .Y(\wave_gen_inst/rom/_193_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_275_  (.A(\wave_gen_inst/rom/_192_ ),
    .B(\wave_gen_inst/rom/_193_ ),
    .Y(\wave_gen_inst/rom/_194_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_276_  (.A(\wave_gen_inst/sine_phase[6] ),
    .B(\wave_gen_inst/rom/_189_ ),
    .C(\wave_gen_inst/rom/_194_ ),
    .Y(\wave_gen_inst/rom/_195_ ));
 sky130_fd_sc_hd__inv_6 \wave_gen_inst/rom/_277_  (.A(\wave_gen_inst/sine_phase[3] ),
    .Y(\wave_gen_inst/rom/_196_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_4 \wave_gen_inst/rom/_279_  (.A(\wave_gen_inst/sine_phase[2] ),
    .SLEEP(\wave_gen_inst/sine_phase[0] ),
    .X(\wave_gen_inst/rom/_198_ ));
 sky130_fd_sc_hd__and2_2 \wave_gen_inst/rom/_280_  (.A(\wave_gen_inst/sine_phase[2] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_199_ ));
 sky130_fd_sc_hd__nand2b_4 \wave_gen_inst/rom/_281_  (.A_N(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_200_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_282_  (.A1(\wave_gen_inst/rom/_198_ ),
    .A2(\wave_gen_inst/rom/_199_ ),
    .B1(\wave_gen_inst/rom/_200_ ),
    .Y(\wave_gen_inst/rom/_201_ ));
 sky130_fd_sc_hd__xor2_1 \wave_gen_inst/rom/_284_  (.A(net71),
    .B(\wave_gen_inst/sine_phase[0] ),
    .X(\wave_gen_inst/rom/_203_ ));
 sky130_fd_sc_hd__o221ai_1 \wave_gen_inst/rom/_286_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/rom/_201_ ),
    .B1(\wave_gen_inst/rom/_203_ ),
    .B2(\wave_gen_inst/sine_phase[2] ),
    .C1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_205_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/rom/_288_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_207_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_289_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/rom/_200_ ),
    .B1(\wave_gen_inst/rom/_207_ ),
    .Y(\wave_gen_inst/rom/_208_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_290_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_209_ ));
 sky130_fd_sc_hd__o31a_1 \wave_gen_inst/rom/_291_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[2] ),
    .A3(\wave_gen_inst/sine_phase[1] ),
    .B1(\wave_gen_inst/sine_phase[3] ),
    .X(\wave_gen_inst/rom/_210_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_292_  (.A1(\wave_gen_inst/rom/_209_ ),
    .A2(\wave_gen_inst/rom/_210_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_211_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_293_  (.A1(net70),
    .A2(\wave_gen_inst/rom/_208_ ),
    .B1(\wave_gen_inst/rom/_211_ ),
    .Y(\wave_gen_inst/rom/_212_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_295_  (.A1(\wave_gen_inst/rom/_205_ ),
    .A2(\wave_gen_inst/rom/_212_ ),
    .B1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_214_ ));
 sky130_fd_sc_hd__nand2b_2 \wave_gen_inst/rom/_296_  (.A_N(\wave_gen_inst/sine_phase[1] ),
    .B(\wave_gen_inst/sine_phase[0] ),
    .Y(\wave_gen_inst/rom/_215_ ));
 sky130_fd_sc_hd__nand4_4 \wave_gen_inst/rom/_297_  (.A(\wave_gen_inst/rom/_196_ ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/rom/_215_ ),
    .D(\wave_gen_inst/rom/_200_ ),
    .Y(\wave_gen_inst/rom/_216_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_299_  (.A(net71),
    .B(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_218_ ));
 sky130_fd_sc_hd__a21bo_1 \wave_gen_inst/rom/_300_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1_N(net71),
    .X(\wave_gen_inst/rom/_219_ ));
 sky130_fd_sc_hd__or2_1 \wave_gen_inst/rom/_301_  (.A(\wave_gen_inst/rom/_198_ ),
    .B(\wave_gen_inst/rom/_219_ ),
    .X(\wave_gen_inst/rom/_220_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/rom/_302_  (.A1(\wave_gen_inst/rom/_200_ ),
    .A2(\wave_gen_inst/rom/_218_ ),
    .B1(\wave_gen_inst/rom/_220_ ),
    .X(\wave_gen_inst/rom/_221_ ));
 sky130_fd_sc_hd__inv_2 \wave_gen_inst/rom/_303_  (.A(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_222_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/rom/_305_  (.A(\wave_gen_inst/rom/_222_ ),
    .B(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_224_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_307_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(\wave_gen_inst/rom/_184_ ),
    .Y(\wave_gen_inst/rom/_226_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/rom/_308_  (.A1(\wave_gen_inst/rom/_226_ ),
    .A2(\wave_gen_inst/rom/_192_ ),
    .B1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_227_ ));
 sky130_fd_sc_hd__a32oi_4 \wave_gen_inst/rom/_309_  (.A1(\wave_gen_inst/rom/_216_ ),
    .A2(\wave_gen_inst/rom/_221_ ),
    .A3(\wave_gen_inst/rom/_224_ ),
    .B1(\wave_gen_inst/rom/_227_ ),
    .B2(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_228_ ));
 sky130_fd_sc_hd__o32ai_4 \wave_gen_inst/rom/_310_  (.A1(\wave_gen_inst/sine_phase[5] ),
    .A2(\wave_gen_inst/rom/_182_ ),
    .A3(\wave_gen_inst/rom/_195_ ),
    .B1(\wave_gen_inst/rom/_214_ ),
    .B2(\wave_gen_inst/rom/_228_ ),
    .Y(\wave_gen_inst/rom_output[0] ));
 sky130_fd_sc_hd__a21oi_4 \wave_gen_inst/rom/_311_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_229_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_312_  (.A(\wave_gen_inst/rom/_196_ ),
    .B(\wave_gen_inst/rom/_229_ ),
    .Y(\wave_gen_inst/rom/_230_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_313_  (.A(net70),
    .B(\wave_gen_inst/rom/_200_ ),
    .Y(\wave_gen_inst/rom/_231_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/rom/_314_  (.A(\wave_gen_inst/sine_phase[1] ),
    .SLEEP(\wave_gen_inst/sine_phase[0] ),
    .X(\wave_gen_inst/rom/_232_ ));
 sky130_fd_sc_hd__o31ai_2 \wave_gen_inst/rom/_315_  (.A1(\wave_gen_inst/rom/_232_ ),
    .A2(\wave_gen_inst/rom/_198_ ),
    .A3(\wave_gen_inst/rom/_199_ ),
    .B1(net71),
    .Y(\wave_gen_inst/rom/_233_ ));
 sky130_fd_sc_hd__or2_1 \wave_gen_inst/rom/_316_  (.A(net71),
    .B(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_234_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/rom/_317_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/rom/_234_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .X(\wave_gen_inst/rom/_235_ ));
 sky130_fd_sc_hd__a32oi_2 \wave_gen_inst/rom/_318_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_230_ ),
    .A3(\wave_gen_inst/rom/_231_ ),
    .B1(\wave_gen_inst/rom/_233_ ),
    .B2(\wave_gen_inst/rom/_235_ ),
    .Y(\wave_gen_inst/rom/_236_ ));
 sky130_fd_sc_hd__or2_2 \wave_gen_inst/rom/_319_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_237_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_320_  (.A1(\wave_gen_inst/rom/_237_ ),
    .A2(\wave_gen_inst/rom/_229_ ),
    .B1(\wave_gen_inst/rom/_199_ ),
    .Y(\wave_gen_inst/rom/_000_ ));
 sky130_fd_sc_hd__or2_1 \wave_gen_inst/rom/_321_  (.A(\wave_gen_inst/sine_phase[2] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_001_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_322_  (.A(net70),
    .B(\wave_gen_inst/rom/_190_ ),
    .C(\wave_gen_inst/rom/_001_ ),
    .Y(\wave_gen_inst/rom/_002_ ));
 sky130_fd_sc_hd__o211a_1 \wave_gen_inst/rom/_323_  (.A1(net71),
    .A2(\wave_gen_inst/rom/_000_ ),
    .B1(\wave_gen_inst/rom/_002_ ),
    .C1(\wave_gen_inst/sine_phase[4] ),
    .X(\wave_gen_inst/rom/_003_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \wave_gen_inst/rom/_324_  (.A(\wave_gen_inst/sine_phase[2] ),
    .SLEEP(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_004_ ));
 sky130_fd_sc_hd__and2_1 \wave_gen_inst/rom/_325_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .X(\wave_gen_inst/rom/_005_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_2 \wave_gen_inst/rom/_326_  (.A(\wave_gen_inst/sine_phase[1] ),
    .SLEEP(\wave_gen_inst/sine_phase[2] ),
    .X(\wave_gen_inst/rom/_006_ ));
 sky130_fd_sc_hd__o41a_1 \wave_gen_inst/rom/_327_  (.A1(\wave_gen_inst/rom/_004_ ),
    .A2(\wave_gen_inst/rom/_005_ ),
    .A3(\wave_gen_inst/rom/_207_ ),
    .A4(\wave_gen_inst/rom/_006_ ),
    .B1(\wave_gen_inst/sine_phase[3] ),
    .X(\wave_gen_inst/rom/_007_ ));
 sky130_fd_sc_hd__nand2b_4 \wave_gen_inst/rom/_328_  (.A_N(\wave_gen_inst/sine_phase[2] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_008_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_329_  (.A1(\wave_gen_inst/rom/_166_ ),
    .A2(\wave_gen_inst/rom/_008_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_009_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_331_  (.A1(\wave_gen_inst/rom/_007_ ),
    .A2(\wave_gen_inst/rom/_009_ ),
    .B1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_011_ ));
 sky130_fd_sc_hd__o22ai_2 \wave_gen_inst/rom/_332_  (.A1(net68),
    .A2(\wave_gen_inst/rom/_236_ ),
    .B1(\wave_gen_inst/rom/_003_ ),
    .B2(\wave_gen_inst/rom/_011_ ),
    .Y(\wave_gen_inst/rom/_012_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/rom/_333_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/sine_phase[0] ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_013_ ));
 sky130_fd_sc_hd__xnor2_4 \wave_gen_inst/rom/_334_  (.A(\wave_gen_inst/sine_phase[2] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_014_ ));
 sky130_fd_sc_hd__a211o_1 \wave_gen_inst/rom/_335_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/rom/_014_ ),
    .B1(\wave_gen_inst/rom/_232_ ),
    .C1(\wave_gen_inst/rom/_196_ ),
    .X(\wave_gen_inst/rom/_015_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_336_  (.A(net70),
    .B(\wave_gen_inst/rom/_169_ ),
    .Y(\wave_gen_inst/rom/_016_ ));
 sky130_fd_sc_hd__and3_1 \wave_gen_inst/rom/_337_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_017_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_338_  (.A(net70),
    .B(\wave_gen_inst/rom/_207_ ),
    .C(\wave_gen_inst/rom/_017_ ),
    .Y(\wave_gen_inst/rom/_018_ ));
 sky130_fd_sc_hd__o21bai_1 \wave_gen_inst/rom/_339_  (.A1(\wave_gen_inst/sine_phase[1] ),
    .A2(\wave_gen_inst/rom/_016_ ),
    .B1_N(\wave_gen_inst/rom/_018_ ),
    .Y(\wave_gen_inst/rom/_019_ ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/rom/_341_  (.A1(\wave_gen_inst/rom/_013_ ),
    .A2(\wave_gen_inst/rom/_015_ ),
    .B1(\wave_gen_inst/rom/_019_ ),
    .B2(\wave_gen_inst/sine_phase[4] ),
    .C1(net68),
    .X(\wave_gen_inst/rom/_021_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_342_  (.A(net71),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_022_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_343_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_023_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_344_  (.A(net71),
    .B(\wave_gen_inst/rom/_023_ ),
    .Y(\wave_gen_inst/rom/_024_ ));
 sky130_fd_sc_hd__nand4_1 \wave_gen_inst/rom/_345_  (.A(\wave_gen_inst/rom/_234_ ),
    .B(\wave_gen_inst/rom/_013_ ),
    .C(\wave_gen_inst/rom/_022_ ),
    .D(\wave_gen_inst/rom/_024_ ),
    .Y(\wave_gen_inst/rom/_025_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_346_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/rom/_234_ ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_026_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/rom/_347_  (.A1(net71),
    .A2(\wave_gen_inst/sine_phase[0] ),
    .B1(\wave_gen_inst/rom/_175_ ),
    .B2(\wave_gen_inst/rom/_184_ ),
    .Y(\wave_gen_inst/rom/_027_ ));
 sky130_fd_sc_hd__o21a_1 \wave_gen_inst/rom/_349_  (.A1(\wave_gen_inst/rom/_026_ ),
    .A2(\wave_gen_inst/rom/_027_ ),
    .B1(net68),
    .X(\wave_gen_inst/rom/_029_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_350_  (.A1(\wave_gen_inst/rom/_025_ ),
    .A2(\wave_gen_inst/rom/_029_ ),
    .B1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_030_ ));
 sky130_fd_sc_hd__a22oi_4 \wave_gen_inst/rom/_351_  (.A1(\wave_gen_inst/sine_phase[6] ),
    .A2(\wave_gen_inst/rom/_012_ ),
    .B1(\wave_gen_inst/rom/_021_ ),
    .B2(\wave_gen_inst/rom/_030_ ),
    .Y(\wave_gen_inst/rom_output[1] ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_352_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/rom/_014_ ),
    .B1(\wave_gen_inst/rom/_196_ ),
    .Y(\wave_gen_inst/rom/_031_ ));
 sky130_fd_sc_hd__a21boi_1 \wave_gen_inst/rom/_353_  (.A1(\wave_gen_inst/rom/_190_ ),
    .A2(\wave_gen_inst/rom/_191_ ),
    .B1_N(\wave_gen_inst/rom/_215_ ),
    .Y(\wave_gen_inst/rom/_032_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_354_  (.A(\wave_gen_inst/rom/_207_ ),
    .B(\wave_gen_inst/rom/_185_ ),
    .Y(\wave_gen_inst/rom/_033_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/rom/_355_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/rom/_032_ ),
    .B1(\wave_gen_inst/rom/_033_ ),
    .C1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_034_ ));
 sky130_fd_sc_hd__o311a_1 \wave_gen_inst/rom/_356_  (.A1(\wave_gen_inst/sine_phase[5] ),
    .A2(\wave_gen_inst/rom/_031_ ),
    .A3(\wave_gen_inst/rom/_018_ ),
    .B1(\wave_gen_inst/rom/_034_ ),
    .C1(\wave_gen_inst/sine_phase[4] ),
    .X(\wave_gen_inst/rom/_035_ ));
 sky130_fd_sc_hd__xor3_1 \wave_gen_inst/rom/_357_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/sine_phase[1] ),
    .X(\wave_gen_inst/rom/_036_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/rom/_358_  (.A(\wave_gen_inst/sine_phase[3] ),
    .B(\wave_gen_inst/rom/_036_ ),
    .Y(\wave_gen_inst/rom/_037_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_359_  (.A(\wave_gen_inst/sine_phase[3] ),
    .B(\wave_gen_inst/sine_phase[0] ),
    .C(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_038_ ));
 sky130_fd_sc_hd__and3b_1 \wave_gen_inst/rom/_360_  (.A_N(\wave_gen_inst/sine_phase[1] ),
    .B(\wave_gen_inst/sine_phase[2] ),
    .C(\wave_gen_inst/sine_phase[0] ),
    .X(\wave_gen_inst/rom/_039_ ));
 sky130_fd_sc_hd__a2111oi_0 \wave_gen_inst/rom/_361_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(\wave_gen_inst/rom/_207_ ),
    .C1(\wave_gen_inst/rom/_039_ ),
    .D1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_040_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_362_  (.A1(\wave_gen_inst/rom/_038_ ),
    .A2(\wave_gen_inst/rom/_040_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_041_ ));
 sky130_fd_sc_hd__o311ai_2 \wave_gen_inst/rom/_363_  (.A1(\wave_gen_inst/rom/_222_ ),
    .A2(\wave_gen_inst/sine_phase[4] ),
    .A3(\wave_gen_inst/rom/_037_ ),
    .B1(\wave_gen_inst/rom/_041_ ),
    .C1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_042_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_364_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/rom/_014_ ),
    .B1(\wave_gen_inst/sine_phase[3] ),
    .Y(\wave_gen_inst/rom/_043_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_365_  (.A1(\wave_gen_inst/rom/_210_ ),
    .A2(\wave_gen_inst/rom/_185_ ),
    .B1(\wave_gen_inst/rom/_222_ ),
    .Y(\wave_gen_inst/rom/_044_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/rom/_366_  (.A1(\wave_gen_inst/rom/_222_ ),
    .A2(\wave_gen_inst/rom/_007_ ),
    .A3(\wave_gen_inst/rom/_043_ ),
    .B1(\wave_gen_inst/rom/_044_ ),
    .Y(\wave_gen_inst/rom/_045_ ));
 sky130_fd_sc_hd__nor2_2 \wave_gen_inst/rom/_367_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/sine_phase[1] ),
    .Y(\wave_gen_inst/rom/_046_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/rom/_368_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(\wave_gen_inst/sine_phase[2] ),
    .X(\wave_gen_inst/rom/_047_ ));
 sky130_fd_sc_hd__o2111ai_2 \wave_gen_inst/rom/_369_  (.A1(\wave_gen_inst/rom/_046_ ),
    .A2(\wave_gen_inst/rom/_047_ ),
    .B1(\wave_gen_inst/rom/_196_ ),
    .C1(\wave_gen_inst/rom/_191_ ),
    .D1(\wave_gen_inst/rom/_175_ ),
    .Y(\wave_gen_inst/rom/_048_ ));
 sky130_fd_sc_hd__nand2_2 \wave_gen_inst/rom/_370_  (.A(\wave_gen_inst/sine_phase[5] ),
    .B(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_049_ ));
 sky130_fd_sc_hd__o311ai_1 \wave_gen_inst/rom/_371_  (.A1(\wave_gen_inst/sine_phase[3] ),
    .A2(\wave_gen_inst/rom/_039_ ),
    .A3(\wave_gen_inst/rom/_006_ ),
    .B1(\wave_gen_inst/rom/_179_ ),
    .C1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_050_ ));
 sky130_fd_sc_hd__a32oi_1 \wave_gen_inst/rom/_372_  (.A1(\wave_gen_inst/sine_phase[5] ),
    .A2(\wave_gen_inst/rom/_220_ ),
    .A3(\wave_gen_inst/rom/_048_ ),
    .B1(\wave_gen_inst/rom/_049_ ),
    .B2(\wave_gen_inst/rom/_050_ ),
    .Y(\wave_gen_inst/rom/_051_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_373_  (.A1(\wave_gen_inst/rom/_187_ ),
    .A2(\wave_gen_inst/rom/_045_ ),
    .B1(\wave_gen_inst/rom/_051_ ),
    .Y(\wave_gen_inst/rom/_052_ ));
 sky130_fd_sc_hd__o22a_4 \wave_gen_inst/rom/_374_  (.A1(\wave_gen_inst/rom/_035_ ),
    .A2(\wave_gen_inst/rom/_042_ ),
    .B1(\wave_gen_inst/rom/_052_ ),
    .B2(\wave_gen_inst/sine_phase[6] ),
    .X(\wave_gen_inst/rom_output[2] ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_375_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/rom/_200_ ),
    .B1(net71),
    .Y(\wave_gen_inst/rom/_053_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_376_  (.A(\wave_gen_inst/rom/_006_ ),
    .B(\wave_gen_inst/rom/_220_ ),
    .Y(\wave_gen_inst/rom/_054_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/rom/_377_  (.A1(\wave_gen_inst/rom/_237_ ),
    .A2(\wave_gen_inst/rom/_229_ ),
    .B1(\wave_gen_inst/rom/_198_ ),
    .Y(\wave_gen_inst/rom/_055_ ));
 sky130_fd_sc_hd__o31ai_2 \wave_gen_inst/rom/_378_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[2] ),
    .A3(\wave_gen_inst/sine_phase[1] ),
    .B1(net70),
    .Y(\wave_gen_inst/rom/_056_ ));
 sky130_fd_sc_hd__o211ai_4 \wave_gen_inst/rom/_379_  (.A1(net70),
    .A2(\wave_gen_inst/rom/_055_ ),
    .B1(\wave_gen_inst/rom/_056_ ),
    .C1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_057_ ));
 sky130_fd_sc_hd__o311ai_4 \wave_gen_inst/rom/_380_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_053_ ),
    .A3(\wave_gen_inst/rom/_054_ ),
    .B1(\wave_gen_inst/rom/_057_ ),
    .C1(\wave_gen_inst/rom/_222_ ),
    .Y(\wave_gen_inst/rom/_058_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_381_  (.A(\wave_gen_inst/rom/_196_ ),
    .B(\wave_gen_inst/rom/_008_ ),
    .Y(\wave_gen_inst/rom/_059_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/rom/_382_  (.A1(\wave_gen_inst/rom/_059_ ),
    .A2(\wave_gen_inst/rom/_231_ ),
    .B1(\wave_gen_inst/rom/_005_ ),
    .X(\wave_gen_inst/rom/_060_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/rom/_383_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(\wave_gen_inst/sine_phase[2] ),
    .Y(\wave_gen_inst/rom/_061_ ));
 sky130_fd_sc_hd__a22oi_1 \wave_gen_inst/rom/_384_  (.A1(\wave_gen_inst/rom/_207_ ),
    .A2(\wave_gen_inst/rom/_185_ ),
    .B1(\wave_gen_inst/rom/_061_ ),
    .B2(net70),
    .Y(\wave_gen_inst/rom/_062_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_385_  (.A(\wave_gen_inst/rom/_049_ ),
    .B(\wave_gen_inst/rom/_062_ ),
    .Y(\wave_gen_inst/rom/_063_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_386_  (.A1(\wave_gen_inst/rom/_224_ ),
    .A2(\wave_gen_inst/rom/_060_ ),
    .B1(\wave_gen_inst/rom/_063_ ),
    .Y(\wave_gen_inst/rom/_064_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_387_  (.A(\wave_gen_inst/sine_phase[2] ),
    .B(\wave_gen_inst/rom/_200_ ),
    .C(\wave_gen_inst/rom/_219_ ),
    .Y(\wave_gen_inst/rom/_065_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_388_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/rom/_219_ ),
    .B1(\wave_gen_inst/rom/_065_ ),
    .Y(\wave_gen_inst/rom/_066_ ));
 sky130_fd_sc_hd__lpflow_isobufsrc_1 \wave_gen_inst/rom/_389_  (.A(\wave_gen_inst/sine_phase[2] ),
    .SLEEP(net71),
    .X(\wave_gen_inst/rom/_067_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_390_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(\wave_gen_inst/rom/_067_ ),
    .Y(\wave_gen_inst/rom/_068_ ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/rom/_391_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_066_ ),
    .B1(\wave_gen_inst/rom/_068_ ),
    .B2(\wave_gen_inst/rom/_024_ ),
    .C1(\wave_gen_inst/sine_phase[5] ),
    .X(\wave_gen_inst/rom/_069_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_392_  (.A1(net71),
    .A2(\wave_gen_inst/rom/_023_ ),
    .B1(\wave_gen_inst/rom/_233_ ),
    .Y(\wave_gen_inst/rom/_070_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_393_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(net70),
    .Y(\wave_gen_inst/rom/_071_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_394_  (.A(\wave_gen_inst/rom/_219_ ),
    .B(\wave_gen_inst/rom/_169_ ),
    .Y(\wave_gen_inst/rom/_072_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_395_  (.A(\wave_gen_inst/rom/_071_ ),
    .B(\wave_gen_inst/rom/_049_ ),
    .C(\wave_gen_inst/rom/_072_ ),
    .Y(\wave_gen_inst/rom/_073_ ));
 sky130_fd_sc_hd__a211oi_2 \wave_gen_inst/rom/_396_  (.A1(\wave_gen_inst/rom/_224_ ),
    .A2(\wave_gen_inst/rom/_070_ ),
    .B1(\wave_gen_inst/rom/_073_ ),
    .C1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_074_ ));
 sky130_fd_sc_hd__a32oi_4 \wave_gen_inst/rom/_397_  (.A1(\wave_gen_inst/sine_phase[6] ),
    .A2(\wave_gen_inst/rom/_058_ ),
    .A3(\wave_gen_inst/rom/_064_ ),
    .B1(\wave_gen_inst/rom/_069_ ),
    .B2(\wave_gen_inst/rom/_074_ ),
    .Y(\wave_gen_inst/rom_output[3] ));
 sky130_fd_sc_hd__clkinv_4 \wave_gen_inst/rom/_398_  (.A(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_075_ ));
 sky130_fd_sc_hd__nor2b_1 \wave_gen_inst/rom/_399_  (.A(\wave_gen_inst/rom/_193_ ),
    .B_N(\wave_gen_inst/rom/_055_ ),
    .Y(\wave_gen_inst/rom/_076_ ));
 sky130_fd_sc_hd__a21o_1 \wave_gen_inst/rom/_400_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(net70),
    .X(\wave_gen_inst/rom/_077_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_401_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(\wave_gen_inst/rom/_001_ ),
    .Y(\wave_gen_inst/rom/_078_ ));
 sky130_fd_sc_hd__a21o_2 \wave_gen_inst/rom/_402_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(net71),
    .X(\wave_gen_inst/rom/_079_ ));
 sky130_fd_sc_hd__o32ai_4 \wave_gen_inst/rom/_403_  (.A1(\wave_gen_inst/rom/_046_ ),
    .A2(\wave_gen_inst/rom/_077_ ),
    .A3(\wave_gen_inst/rom/_078_ ),
    .B1(\wave_gen_inst/rom/_079_ ),
    .B2(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_080_ ));
 sky130_fd_sc_hd__a31oi_4 \wave_gen_inst/rom/_404_  (.A1(\wave_gen_inst/rom/_216_ ),
    .A2(\wave_gen_inst/rom/_008_ ),
    .A3(\wave_gen_inst/rom/_016_ ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_081_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_405_  (.A1(\wave_gen_inst/rom/_203_ ),
    .A2(\wave_gen_inst/rom/_026_ ),
    .B1(net68),
    .Y(\wave_gen_inst/rom/_082_ ));
 sky130_fd_sc_hd__o32ai_4 \wave_gen_inst/rom/_406_  (.A1(net68),
    .A2(\wave_gen_inst/rom/_076_ ),
    .A3(\wave_gen_inst/rom/_080_ ),
    .B1(\wave_gen_inst/rom/_081_ ),
    .B2(\wave_gen_inst/rom/_082_ ),
    .Y(\wave_gen_inst/rom/_083_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_407_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/sine_phase[1] ),
    .B1(net71),
    .Y(\wave_gen_inst/rom/_084_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_408_  (.A(\wave_gen_inst/sine_phase[0] ),
    .B(\wave_gen_inst/rom/_084_ ),
    .Y(\wave_gen_inst/rom/_085_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_409_  (.A1(\wave_gen_inst/rom/_046_ ),
    .A2(\wave_gen_inst/rom/_047_ ),
    .B1(net70),
    .Y(\wave_gen_inst/rom/_086_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_410_  (.A1(\wave_gen_inst/rom/_085_ ),
    .A2(\wave_gen_inst/rom/_086_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_087_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_411_  (.A(\wave_gen_inst/sine_phase[1] ),
    .B(\wave_gen_inst/rom/_175_ ),
    .Y(\wave_gen_inst/rom/_088_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_412_  (.A1(\wave_gen_inst/rom/_088_ ),
    .A2(\wave_gen_inst/rom/_193_ ),
    .B1(net68),
    .Y(\wave_gen_inst/rom/_089_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/rom/_413_  (.A1(\wave_gen_inst/rom/_209_ ),
    .A2(\wave_gen_inst/rom/_008_ ),
    .A3(\wave_gen_inst/rom/_234_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_090_ ));
 sky130_fd_sc_hd__a22oi_2 \wave_gen_inst/rom/_414_  (.A1(\wave_gen_inst/rom/_002_ ),
    .A2(\wave_gen_inst/rom/_013_ ),
    .B1(\wave_gen_inst/rom/_085_ ),
    .B2(\wave_gen_inst/rom/_090_ ),
    .Y(\wave_gen_inst/rom/_091_ ));
 sky130_fd_sc_hd__o221ai_4 \wave_gen_inst/rom/_415_  (.A1(\wave_gen_inst/rom/_087_ ),
    .A2(\wave_gen_inst/rom/_089_ ),
    .B1(\wave_gen_inst/rom/_091_ ),
    .B2(net68),
    .C1(\wave_gen_inst/rom/_075_ ),
    .Y(\wave_gen_inst/rom/_092_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/rom/_416_  (.A1(\wave_gen_inst/rom/_075_ ),
    .A2(\wave_gen_inst/rom/_083_ ),
    .B1(\wave_gen_inst/rom/_092_ ),
    .Y(\wave_gen_inst/rom_output[4] ));
 sky130_fd_sc_hd__a221o_1 \wave_gen_inst/rom/_417_  (.A1(\wave_gen_inst/sine_phase[2] ),
    .A2(\wave_gen_inst/rom/_215_ ),
    .B1(\wave_gen_inst/rom/_237_ ),
    .B2(\wave_gen_inst/rom/_229_ ),
    .C1(net70),
    .X(\wave_gen_inst/rom/_093_ ));
 sky130_fd_sc_hd__o211a_1 \wave_gen_inst/rom/_418_  (.A1(\wave_gen_inst/rom/_004_ ),
    .A2(\wave_gen_inst/rom/_086_ ),
    .B1(\wave_gen_inst/rom/_093_ ),
    .C1(\wave_gen_inst/rom/_187_ ),
    .X(\wave_gen_inst/rom/_094_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_419_  (.A1(\wave_gen_inst/rom/_046_ ),
    .A2(\wave_gen_inst/rom/_077_ ),
    .B1(\wave_gen_inst/rom/_184_ ),
    .Y(\wave_gen_inst/rom/_095_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_420_  (.A1(\wave_gen_inst/rom/_187_ ),
    .A2(\wave_gen_inst/rom/_095_ ),
    .B1(net68),
    .Y(\wave_gen_inst/rom/_097_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/rom/_421_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/rom/_014_ ),
    .B1(\wave_gen_inst/rom/_198_ ),
    .C1(\wave_gen_inst/sine_phase[3] ),
    .Y(\wave_gen_inst/rom/_098_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_422_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/sine_phase[0] ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_099_ ));
 sky130_fd_sc_hd__o32ai_2 \wave_gen_inst/rom/_423_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_196_ ),
    .A3(\wave_gen_inst/rom/_032_ ),
    .B1(\wave_gen_inst/rom/_098_ ),
    .B2(\wave_gen_inst/rom/_099_ ),
    .Y(\wave_gen_inst/rom/_100_ ));
 sky130_fd_sc_hd__o22ai_1 \wave_gen_inst/rom/_424_  (.A1(\wave_gen_inst/rom/_094_ ),
    .A2(\wave_gen_inst/rom/_097_ ),
    .B1(\wave_gen_inst/rom/_100_ ),
    .B2(net68),
    .Y(\wave_gen_inst/rom/_101_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_425_  (.A1(\wave_gen_inst/rom/_210_ ),
    .A2(\wave_gen_inst/rom/_185_ ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_102_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_426_  (.A(\wave_gen_inst/rom/_013_ ),
    .B(\wave_gen_inst/rom/_037_ ),
    .Y(\wave_gen_inst/rom/_103_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_427_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(net70),
    .Y(\wave_gen_inst/rom/_104_ ));
 sky130_fd_sc_hd__a2111oi_0 \wave_gen_inst/rom/_428_  (.A1(\wave_gen_inst/rom/_237_ ),
    .A2(\wave_gen_inst/rom/_229_ ),
    .B1(\wave_gen_inst/rom/_104_ ),
    .C1(\wave_gen_inst/rom/_199_ ),
    .D1(\wave_gen_inst/rom/_198_ ),
    .Y(\wave_gen_inst/rom/_105_ ));
 sky130_fd_sc_hd__nor4_1 \wave_gen_inst/rom/_429_  (.A(\wave_gen_inst/rom/_187_ ),
    .B(\wave_gen_inst/rom/_198_ ),
    .C(\wave_gen_inst/rom/_046_ ),
    .D(\wave_gen_inst/rom/_077_ ),
    .Y(\wave_gen_inst/rom/_106_ ));
 sky130_fd_sc_hd__a2111oi_0 \wave_gen_inst/rom/_430_  (.A1(\wave_gen_inst/rom/_187_ ),
    .A2(\wave_gen_inst/rom/_095_ ),
    .B1(\wave_gen_inst/rom/_105_ ),
    .C1(\wave_gen_inst/rom/_106_ ),
    .D1(net68),
    .Y(\wave_gen_inst/rom/_108_ ));
 sky130_fd_sc_hd__a311oi_1 \wave_gen_inst/rom/_431_  (.A1(net68),
    .A2(\wave_gen_inst/rom/_102_ ),
    .A3(\wave_gen_inst/rom/_103_ ),
    .B1(\wave_gen_inst/rom/_108_ ),
    .C1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_109_ ));
 sky130_fd_sc_hd__a21o_4 \wave_gen_inst/rom/_432_  (.A1(\wave_gen_inst/sine_phase[6] ),
    .A2(\wave_gen_inst/rom/_101_ ),
    .B1(\wave_gen_inst/rom/_109_ ),
    .X(\wave_gen_inst/rom_output[5] ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_433_  (.A1(\wave_gen_inst/rom/_001_ ),
    .A2(\wave_gen_inst/rom/_061_ ),
    .B1(net70),
    .Y(\wave_gen_inst/rom/_110_ ));
 sky130_fd_sc_hd__o32a_1 \wave_gen_inst/rom/_434_  (.A1(\wave_gen_inst/rom/_193_ ),
    .A2(\wave_gen_inst/rom/_229_ ),
    .A3(\wave_gen_inst/rom/_017_ ),
    .B1(\wave_gen_inst/rom/_110_ ),
    .B2(\wave_gen_inst/rom/_226_ ),
    .X(\wave_gen_inst/rom/_111_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_435_  (.A(\wave_gen_inst/rom/_075_ ),
    .B(\wave_gen_inst/rom/_111_ ),
    .Y(\wave_gen_inst/rom/_112_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_436_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(\wave_gen_inst/rom/_037_ ),
    .Y(\wave_gen_inst/rom/_113_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_437_  (.A1(\wave_gen_inst/rom/_192_ ),
    .A2(\wave_gen_inst/rom/_008_ ),
    .B1(\wave_gen_inst/rom/_104_ ),
    .Y(\wave_gen_inst/rom/_114_ ));
 sky130_fd_sc_hd__a211oi_1 \wave_gen_inst/rom/_438_  (.A1(\wave_gen_inst/rom/_190_ ),
    .A2(\wave_gen_inst/rom/_006_ ),
    .B1(\wave_gen_inst/rom/_005_ ),
    .C1(\wave_gen_inst/rom/_004_ ),
    .Y(\wave_gen_inst/rom/_115_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_439_  (.A1(net70),
    .A2(\wave_gen_inst/rom/_115_ ),
    .B1(\wave_gen_inst/rom/_075_ ),
    .Y(\wave_gen_inst/rom/_116_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_440_  (.A(\wave_gen_inst/rom/_113_ ),
    .B(\wave_gen_inst/rom/_114_ ),
    .C(\wave_gen_inst/rom/_116_ ),
    .Y(\wave_gen_inst/rom/_118_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_441_  (.A1(\wave_gen_inst/sine_phase[3] ),
    .A2(\wave_gen_inst/rom/_169_ ),
    .B1(\wave_gen_inst/rom/_098_ ),
    .Y(\wave_gen_inst/rom/_119_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_442_  (.A(\wave_gen_inst/rom/_237_ ),
    .B(\wave_gen_inst/rom/_001_ ),
    .C(\wave_gen_inst/rom/_071_ ),
    .Y(\wave_gen_inst/rom/_120_ ));
 sky130_fd_sc_hd__o211ai_1 \wave_gen_inst/rom/_443_  (.A1(\wave_gen_inst/sine_phase[0] ),
    .A2(\wave_gen_inst/rom/_008_ ),
    .B1(\wave_gen_inst/rom/_175_ ),
    .C1(net70),
    .Y(\wave_gen_inst/rom/_121_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_444_  (.A1(\wave_gen_inst/rom/_120_ ),
    .A2(\wave_gen_inst/rom/_121_ ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_122_ ));
 sky130_fd_sc_hd__a211oi_2 \wave_gen_inst/rom/_445_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_119_ ),
    .B1(\wave_gen_inst/rom/_122_ ),
    .C1(\wave_gen_inst/rom/_075_ ),
    .Y(\wave_gen_inst/rom/_123_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_446_  (.A(\wave_gen_inst/rom/_046_ ),
    .B(\wave_gen_inst/rom/_077_ ),
    .Y(\wave_gen_inst/rom/_124_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_447_  (.A(\wave_gen_inst/rom/_004_ ),
    .B(\wave_gen_inst/rom/_198_ ),
    .C(\wave_gen_inst/rom/_056_ ),
    .Y(\wave_gen_inst/rom/_125_ ));
 sky130_fd_sc_hd__o32a_1 \wave_gen_inst/rom/_448_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_124_ ),
    .A3(\wave_gen_inst/rom/_125_ ),
    .B1(\wave_gen_inst/rom/_079_ ),
    .B2(\wave_gen_inst/rom/_078_ ),
    .X(\wave_gen_inst/rom/_126_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_449_  (.A1(\wave_gen_inst/sine_phase[6] ),
    .A2(\wave_gen_inst/rom/_126_ ),
    .B1(net68),
    .Y(\wave_gen_inst/rom/_127_ ));
 sky130_fd_sc_hd__o32ai_4 \wave_gen_inst/rom/_450_  (.A1(net68),
    .A2(\wave_gen_inst/rom/_112_ ),
    .A3(\wave_gen_inst/rom/_118_ ),
    .B1(\wave_gen_inst/rom/_123_ ),
    .B2(\wave_gen_inst/rom/_127_ ),
    .Y(\wave_gen_inst/rom_output[6] ));
 sky130_fd_sc_hd__or3_1 \wave_gen_inst/rom/_451_  (.A(net71),
    .B(\wave_gen_inst/rom/_004_ ),
    .C(\wave_gen_inst/rom/_023_ ),
    .X(\wave_gen_inst/rom/_129_ ));
 sky130_fd_sc_hd__a221oi_1 \wave_gen_inst/rom/_452_  (.A1(\wave_gen_inst/rom/_067_ ),
    .A2(\wave_gen_inst/rom/_237_ ),
    .B1(\wave_gen_inst/rom/_014_ ),
    .B2(net71),
    .C1(net68),
    .Y(\wave_gen_inst/rom/_130_ ));
 sky130_fd_sc_hd__a31oi_2 \wave_gen_inst/rom/_453_  (.A1(net68),
    .A2(\wave_gen_inst/rom/_015_ ),
    .A3(\wave_gen_inst/rom/_129_ ),
    .B1(\wave_gen_inst/rom/_130_ ),
    .Y(\wave_gen_inst/rom/_131_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_454_  (.A1(\wave_gen_inst/rom/_219_ ),
    .A2(\wave_gen_inst/rom/_229_ ),
    .B1(net68),
    .Y(\wave_gen_inst/rom/_132_ ));
 sky130_fd_sc_hd__o32a_1 \wave_gen_inst/rom/_455_  (.A1(net68),
    .A2(\wave_gen_inst/rom/_175_ ),
    .A3(\wave_gen_inst/rom/_184_ ),
    .B1(\wave_gen_inst/rom/_110_ ),
    .B2(\wave_gen_inst/rom/_132_ ),
    .X(\wave_gen_inst/rom/_133_ ));
 sky130_fd_sc_hd__mux2i_4 \wave_gen_inst/rom/_456_  (.A0(\wave_gen_inst/rom/_131_ ),
    .A1(\wave_gen_inst/rom/_133_ ),
    .S(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_134_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_457_  (.A1(net71),
    .A2(\wave_gen_inst/sine_phase[2] ),
    .B1(\wave_gen_inst/sine_phase[4] ),
    .Y(\wave_gen_inst/rom/_135_ ));
 sky130_fd_sc_hd__o31ai_1 \wave_gen_inst/rom/_458_  (.A1(net71),
    .A2(\wave_gen_inst/rom/_229_ ),
    .A3(\wave_gen_inst/rom/_017_ ),
    .B1(\wave_gen_inst/rom/_135_ ),
    .Y(\wave_gen_inst/rom/_136_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_459_  (.A(net68),
    .B(\wave_gen_inst/rom/_026_ ),
    .C(\wave_gen_inst/rom/_136_ ),
    .Y(\wave_gen_inst/rom/_137_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_460_  (.A1(\wave_gen_inst/rom/_047_ ),
    .A2(\wave_gen_inst/rom/_061_ ),
    .B1(\wave_gen_inst/rom/_193_ ),
    .Y(\wave_gen_inst/rom/_139_ ));
 sky130_fd_sc_hd__nor3_1 \wave_gen_inst/rom/_461_  (.A(net70),
    .B(\wave_gen_inst/rom/_207_ ),
    .C(\wave_gen_inst/rom/_014_ ),
    .Y(\wave_gen_inst/rom/_140_ ));
 sky130_fd_sc_hd__a2111o_1 \wave_gen_inst/rom/_462_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_125_ ),
    .B1(\wave_gen_inst/rom/_139_ ),
    .C1(\wave_gen_inst/rom/_140_ ),
    .D1(net68),
    .X(\wave_gen_inst/rom/_141_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_463_  (.A1(\wave_gen_inst/rom/_137_ ),
    .A2(\wave_gen_inst/rom/_141_ ),
    .B1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_142_ ));
 sky130_fd_sc_hd__a21oi_4 \wave_gen_inst/rom/_464_  (.A1(\wave_gen_inst/sine_phase[6] ),
    .A2(\wave_gen_inst/rom/_134_ ),
    .B1(\wave_gen_inst/rom/_142_ ),
    .Y(\wave_gen_inst/rom_output[7] ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/rom/_465_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/rom/_229_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_143_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_466_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_022_ ),
    .B1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_144_ ));
 sky130_fd_sc_hd__a221oi_2 \wave_gen_inst/rom/_467_  (.A1(\wave_gen_inst/rom/_196_ ),
    .A2(\wave_gen_inst/rom/_061_ ),
    .B1(\wave_gen_inst/rom/_143_ ),
    .B2(\wave_gen_inst/sine_phase[5] ),
    .C1(\wave_gen_inst/rom/_144_ ),
    .Y(\wave_gen_inst/rom/_145_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_468_  (.A(\wave_gen_inst/rom/_196_ ),
    .B(\wave_gen_inst/rom/_229_ ),
    .Y(\wave_gen_inst/rom/_146_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_469_  (.A(\wave_gen_inst/rom/_023_ ),
    .B(\wave_gen_inst/rom/_079_ ),
    .Y(\wave_gen_inst/rom/_147_ ));
 sky130_fd_sc_hd__nor2_1 \wave_gen_inst/rom/_470_  (.A(\wave_gen_inst/rom/_146_ ),
    .B(\wave_gen_inst/rom/_147_ ),
    .Y(\wave_gen_inst/rom/_149_ ));
 sky130_fd_sc_hd__o21ai_2 \wave_gen_inst/rom/_471_  (.A1(\wave_gen_inst/rom/_049_ ),
    .A2(\wave_gen_inst/rom/_149_ ),
    .B1(\wave_gen_inst/sine_phase[6] ),
    .Y(\wave_gen_inst/rom/_150_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_472_  (.A(\wave_gen_inst/sine_phase[4] ),
    .B(\wave_gen_inst/rom/_218_ ),
    .C(\wave_gen_inst/rom/_079_ ),
    .Y(\wave_gen_inst/rom/_151_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_473_  (.A1(\wave_gen_inst/rom/_084_ ),
    .A2(\wave_gen_inst/rom/_146_ ),
    .B1(\wave_gen_inst/rom/_187_ ),
    .Y(\wave_gen_inst/rom/_152_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/rom/_474_  (.A1(\wave_gen_inst/rom/_151_ ),
    .A2(\wave_gen_inst/rom/_152_ ),
    .B1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_153_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_475_  (.A(\wave_gen_inst/rom/_230_ ),
    .B(\wave_gen_inst/rom/_135_ ),
    .Y(\wave_gen_inst/rom/_154_ ));
 sky130_fd_sc_hd__o21ai_1 \wave_gen_inst/rom/_476_  (.A1(\wave_gen_inst/rom/_222_ ),
    .A2(\wave_gen_inst/rom/_154_ ),
    .B1(\wave_gen_inst/rom/_075_ ),
    .Y(\wave_gen_inst/rom/_155_ ));
 sky130_fd_sc_hd__o22ai_4 \wave_gen_inst/rom/_477_  (.A1(\wave_gen_inst/rom/_145_ ),
    .A2(\wave_gen_inst/rom/_150_ ),
    .B1(\wave_gen_inst/rom/_153_ ),
    .B2(\wave_gen_inst/rom/_155_ ),
    .Y(\wave_gen_inst/rom_output[8] ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_478_  (.A(\wave_gen_inst/sine_phase[5] ),
    .B(\wave_gen_inst/rom/_143_ ),
    .Y(\wave_gen_inst/rom/_156_ ));
 sky130_fd_sc_hd__a21oi_1 \wave_gen_inst/rom/_479_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_079_ ),
    .B1(\wave_gen_inst/rom/_156_ ),
    .Y(\wave_gen_inst/rom/_157_ ));
 sky130_fd_sc_hd__a31oi_1 \wave_gen_inst/rom/_480_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(net71),
    .A3(\wave_gen_inst/rom/_199_ ),
    .B1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_159_ ));
 sky130_fd_sc_hd__a21oi_2 \wave_gen_inst/rom/_481_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_079_ ),
    .B1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_160_ ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_482_  (.A(\wave_gen_inst/rom/_143_ ),
    .B(\wave_gen_inst/rom/_160_ ),
    .Y(\wave_gen_inst/rom/_161_ ));
 sky130_fd_sc_hd__o21ai_0 \wave_gen_inst/rom/_483_  (.A1(\wave_gen_inst/sine_phase[4] ),
    .A2(\wave_gen_inst/rom/_230_ ),
    .B1(\wave_gen_inst/sine_phase[5] ),
    .Y(\wave_gen_inst/rom/_162_ ));
 sky130_fd_sc_hd__nand3_1 \wave_gen_inst/rom/_484_  (.A(\wave_gen_inst/rom/_075_ ),
    .B(\wave_gen_inst/rom/_161_ ),
    .C(\wave_gen_inst/rom/_162_ ),
    .Y(\wave_gen_inst/rom/_163_ ));
 sky130_fd_sc_hd__o31a_4 \wave_gen_inst/rom/_485_  (.A1(\wave_gen_inst/rom/_075_ ),
    .A2(\wave_gen_inst/rom/_157_ ),
    .A3(\wave_gen_inst/rom/_159_ ),
    .B1(\wave_gen_inst/rom/_163_ ),
    .X(\wave_gen_inst/rom_output[9] ));
 sky130_fd_sc_hd__nand2_1 \wave_gen_inst/rom/_486_  (.A(\wave_gen_inst/sine_phase[6] ),
    .B(\wave_gen_inst/rom/_156_ ),
    .Y(\wave_gen_inst/rom/_164_ ));
 sky130_fd_sc_hd__o21ai_4 \wave_gen_inst/rom/_487_  (.A1(\wave_gen_inst/sine_phase[6] ),
    .A2(\wave_gen_inst/rom/_160_ ),
    .B1(\wave_gen_inst/rom/_164_ ),
    .Y(\wave_gen_inst/rom_output[10] ));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0743__488  (.A(clknet_leaf_73_clk),
    .Y(net488));
 sky130_fd_sc_hd__buf_1 input1 (.A(ser_rx),
    .X(net1));
 sky130_fd_sc_hd__buf_16 output2 (.A(net2),
    .X(flash_clk));
 sky130_fd_sc_hd__buf_16 output3 (.A(net3),
    .X(flash_csb));
 sky130_fd_sc_hd__buf_16 output4 (.A(net4),
    .X(led1));
 sky130_fd_sc_hd__buf_16 output5 (.A(net5),
    .X(led2));
 sky130_fd_sc_hd__buf_16 output6 (.A(net6),
    .X(led3));
 sky130_fd_sc_hd__buf_16 output7 (.A(net7),
    .X(led4));
 sky130_fd_sc_hd__buf_16 output8 (.A(net8),
    .X(led5));
 sky130_fd_sc_hd__buf_16 output9 (.A(net9),
    .X(ledg_n));
 sky130_fd_sc_hd__buf_16 output10 (.A(net10),
    .X(ledr_n));
 sky130_fd_sc_hd__buf_16 output11 (.A(net11),
    .X(mode[0]));
 sky130_fd_sc_hd__buf_16 output12 (.A(net12),
    .X(mode[1]));
 sky130_fd_sc_hd__buf_16 output13 (.A(net13),
    .X(mode[2]));
 sky130_fd_sc_hd__buf_16 output14 (.A(net14),
    .X(ser_tx));
 sky130_fd_sc_hd__buf_16 output15 (.A(net15),
    .X(wave[0]));
 sky130_fd_sc_hd__buf_16 output16 (.A(net16),
    .X(wave[10]));
 sky130_fd_sc_hd__buf_16 output17 (.A(net17),
    .X(wave[11]));
 sky130_fd_sc_hd__buf_16 output18 (.A(net18),
    .X(wave[12]));
 sky130_fd_sc_hd__buf_16 output19 (.A(net19),
    .X(wave[13]));
 sky130_fd_sc_hd__buf_16 output20 (.A(net20),
    .X(wave[14]));
 sky130_fd_sc_hd__buf_16 output21 (.A(net21),
    .X(wave[15]));
 sky130_fd_sc_hd__buf_16 output22 (.A(net22),
    .X(wave[16]));
 sky130_fd_sc_hd__buf_16 output23 (.A(net23),
    .X(wave[17]));
 sky130_fd_sc_hd__buf_16 output24 (.A(net24),
    .X(wave[18]));
 sky130_fd_sc_hd__buf_16 output25 (.A(net25),
    .X(wave[19]));
 sky130_fd_sc_hd__buf_16 output26 (.A(net26),
    .X(wave[1]));
 sky130_fd_sc_hd__buf_16 output27 (.A(net27),
    .X(wave[20]));
 sky130_fd_sc_hd__buf_16 output28 (.A(net28),
    .X(wave[21]));
 sky130_fd_sc_hd__buf_16 output29 (.A(net29),
    .X(wave[22]));
 sky130_fd_sc_hd__buf_16 output30 (.A(net30),
    .X(wave[23]));
 sky130_fd_sc_hd__buf_16 output31 (.A(net31),
    .X(wave[24]));
 sky130_fd_sc_hd__buf_16 output32 (.A(net32),
    .X(wave[25]));
 sky130_fd_sc_hd__buf_16 output33 (.A(net33),
    .X(wave[26]));
 sky130_fd_sc_hd__buf_16 output34 (.A(net34),
    .X(wave[27]));
 sky130_fd_sc_hd__buf_16 output35 (.A(net35),
    .X(wave[28]));
 sky130_fd_sc_hd__buf_16 output36 (.A(net36),
    .X(wave[29]));
 sky130_fd_sc_hd__buf_16 output37 (.A(net37),
    .X(wave[2]));
 sky130_fd_sc_hd__buf_16 output38 (.A(net38),
    .X(wave[30]));
 sky130_fd_sc_hd__buf_16 output39 (.A(net39),
    .X(wave[31]));
 sky130_fd_sc_hd__buf_16 output40 (.A(net40),
    .X(wave[3]));
 sky130_fd_sc_hd__buf_16 output41 (.A(net41),
    .X(wave[4]));
 sky130_fd_sc_hd__buf_16 output42 (.A(net42),
    .X(wave[5]));
 sky130_fd_sc_hd__buf_16 output43 (.A(net43),
    .X(wave[6]));
 sky130_fd_sc_hd__buf_16 output44 (.A(net44),
    .X(wave[7]));
 sky130_fd_sc_hd__buf_16 output45 (.A(net45),
    .X(wave[8]));
 sky130_fd_sc_hd__buf_16 output46 (.A(net46),
    .X(wave[9]));
 sky130_fd_sc_hd__clkbuf_8 wire47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_8 load_slew48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 wire49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 wire50 (.A(\soc/cpu/_02606_ ),
    .X(net50));
 sky130_fd_sc_hd__buf_8 wire51 (.A(\soc/cpu/_02712_ ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_8 load_slew52 (.A(\soc/cpu/cpuregs_wrdata[29] ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 load_slew53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 load_slew54 (.A(\soc/cpu/_03699_ ),
    .X(net54));
 sky130_fd_sc_hd__buf_6 max_cap55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 wire56 (.A(\soc/cpu/cpuregs_wrdata[27] ),
    .X(net56));
 sky130_fd_sc_hd__buf_6 load_slew57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__buf_8 wire58 (.A(\soc/cpu/cpuregs_wrdata[25] ),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_16 wire59 (.A(\soc/cpu/cpuregs_wrdata[21] ),
    .X(net59));
 sky130_fd_sc_hd__buf_6 max_cap60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 wire61 (.A(\soc/cpu/cpuregs_wrdata[22] ),
    .X(net61));
 sky130_fd_sc_hd__buf_16 max_cap62 (.A(\soc/simpleuart/_0607_ ),
    .X(net62));
 sky130_fd_sc_hd__buf_6 load_slew63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_8 wire64 (.A(\soc/cpu/cpuregs_wrdata[20] ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 load_slew65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_8 load_slew66 (.A(\soc/cpu/_00721_ ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 wire67 (.A(net910),
    .X(net67));
 sky130_fd_sc_hd__buf_6 load_slew68 (.A(\wave_gen_inst/sine_phase[5] ),
    .X(net68));
 sky130_fd_sc_hd__buf_6 load_slew69 (.A(\soc/cpu/cpuregs_wrdata[16] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 load_slew70 (.A(\wave_gen_inst/sine_phase[3] ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 max_cap71 (.A(\wave_gen_inst/sine_phase[3] ),
    .X(net71));
 sky130_fd_sc_hd__buf_12 load_slew72 (.A(\soc/cpu/cpuregs/_2511_ ),
    .X(net72));
 sky130_fd_sc_hd__buf_16 load_slew73 (.A(\soc/cpu/cpuregs/_2511_ ),
    .X(net73));
 sky130_fd_sc_hd__buf_16 load_slew74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_16 max_cap75 (.A(\soc/cpu/cpuregs/_2487_ ),
    .X(net75));
 sky130_fd_sc_hd__buf_16 load_slew76 (.A(\soc/cpu/cpuregs/_2470_ ),
    .X(net76));
 sky130_fd_sc_hd__buf_16 load_slew77 (.A(\soc/cpu/cpuregs/_2470_ ),
    .X(net77));
 sky130_fd_sc_hd__buf_12 load_slew78 (.A(\soc/cpu/cpuregs/_2466_ ),
    .X(net78));
 sky130_fd_sc_hd__buf_12 load_slew79 (.A(\soc/cpu/cpuregs/_2466_ ),
    .X(net79));
 sky130_fd_sc_hd__buf_16 load_slew80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_16 wire81 (.A(\soc/cpu/cpuregs/_2427_ ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_16 load_slew82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_16 load_slew83 (.A(\soc/cpu/cpuregs/_2422_ ),
    .X(net83));
 sky130_fd_sc_hd__buf_16 wire84 (.A(\soc/cpu/cpuregs/_2417_ ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_16 load_slew85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_16 load_slew86 (.A(\soc/cpu/cpuregs/_2373_ ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_8 load_slew87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_8 wire88 (.A(\soc/cpu/cpuregs_wrdata[17] ),
    .X(net88));
 sky130_fd_sc_hd__buf_16 load_slew89 (.A(\soc/cpu/cpuregs/_2495_ ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_16 max_cap90 (.A(\soc/cpu/cpuregs/_2495_ ),
    .X(net90));
 sky130_fd_sc_hd__buf_16 load_slew91 (.A(\soc/cpu/cpuregs/_2474_ ),
    .X(net91));
 sky130_fd_sc_hd__buf_12 load_slew92 (.A(\soc/cpu/cpuregs/_2474_ ),
    .X(net92));
 sky130_fd_sc_hd__buf_16 load_slew93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_12 load_slew94 (.A(\soc/cpu/cpuregs/_2444_ ),
    .X(net94));
 sky130_fd_sc_hd__buf_12 load_slew95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_16 load_slew96 (.A(\soc/cpu/cpuregs/_2440_ ),
    .X(net96));
 sky130_fd_sc_hd__buf_16 load_slew97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__buf_12 load_slew98 (.A(\soc/cpu/cpuregs/_2382_ ),
    .X(net98));
 sky130_fd_sc_hd__buf_12 load_slew99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__buf_12 load_slew100 (.A(\soc/cpu/cpuregs/_2377_ ),
    .X(net100));
 sky130_fd_sc_hd__buf_12 load_slew101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__buf_12 load_slew102 (.A(\soc/cpu/cpuregs/_2362_ ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_16 load_slew103 (.A(\soc/cpu/cpuregs/_2279_ ),
    .X(net103));
 sky130_fd_sc_hd__buf_16 load_slew104 (.A(\soc/cpu/cpuregs/_2279_ ),
    .X(net104));
 sky130_fd_sc_hd__buf_12 wire105 (.A(\soc/cpu/cpuregs_wrdata[13] ),
    .X(net105));
 sky130_fd_sc_hd__buf_12 max_cap106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_16 wire107 (.A(\soc/spimemio/_0305_ ),
    .X(net107));
 sky130_fd_sc_hd__buf_4 load_slew108 (.A(net112),
    .X(net108));
 sky130_fd_sc_hd__buf_4 load_slew109 (.A(net112),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 load_slew110 (.A(\soc/spimem_ready ),
    .X(net110));
 sky130_fd_sc_hd__buf_6 load_slew111 (.A(\soc/spimem_ready ),
    .X(net111));
 sky130_fd_sc_hd__buf_6 max_cap112 (.A(net828),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_8 load_slew113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 wire114 (.A(\soc/cpu/cpuregs_wrdata[14] ),
    .X(net114));
 sky130_fd_sc_hd__buf_2 wire115 (.A(\soc/cpu/_03851_ ),
    .X(net115));
 sky130_fd_sc_hd__buf_2 wire116 (.A(\soc/cpu/_03665_ ),
    .X(net116));
 sky130_fd_sc_hd__buf_2 wire117 (.A(\soc/cpu/_03648_ ),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 wire118 (.A(\soc/cpu/_03634_ ),
    .X(net118));
 sky130_fd_sc_hd__buf_2 wire119 (.A(\soc/cpu/_03603_ ),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_8 wire120 (.A(_088_),
    .X(net120));
 sky130_fd_sc_hd__buf_6 max_cap121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_4 load_slew122 (.A(_088_),
    .X(net122));
 sky130_fd_sc_hd__buf_6 load_slew123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_8 wire124 (.A(\soc/cpu/cpuregs_wrdata[11] ),
    .X(net124));
 sky130_fd_sc_hd__buf_16 wire125 (.A(\soc/cpu/cpuregs_wrdata[7] ),
    .X(net125));
 sky130_fd_sc_hd__buf_6 max_cap126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_8 wire127 (.A(\soc/cpu/cpuregs_wrdata[8] ),
    .X(net127));
 sky130_fd_sc_hd__buf_16 wire128 (.A(\soc/cpu/cpuregs_wrdata[4] ),
    .X(net128));
 sky130_fd_sc_hd__buf_12 wire129 (.A(\soc/cpu/cpuregs_wrdata[3] ),
    .X(net129));
 sky130_fd_sc_hd__buf_16 wire130 (.A(\soc/cpu/cpuregs_wrdata[1] ),
    .X(net130));
 sky130_fd_sc_hd__buf_16 load_slew131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_16 load_slew132 (.A(\soc/cpu/_00840_ ),
    .X(net132));
 sky130_fd_sc_hd__buf_6 max_cap133 (.A(\soc/cpu/_00713_ ),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 wire134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_8 load_slew135 (.A(net742),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_8 load_slew136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_4 load_slew137 (.A(net905),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 load_slew138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_4 load_slew139 (.A(\soc/_025_ ),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 load_slew140 (.A(\wave_gen_inst/_0602_ ),
    .X(net140));
 sky130_fd_sc_hd__buf_4 load_slew141 (.A(\wave_gen_inst/_0602_ ),
    .X(net141));
 sky130_fd_sc_hd__buf_16 max_cap142 (.A(\wave_gen_inst/_0167_ ),
    .X(net142));
 sky130_fd_sc_hd__buf_8 load_slew143 (.A(\soc/cpu/_02554_ ),
    .X(net143));
 sky130_fd_sc_hd__buf_8 load_slew144 (.A(\soc/cpu/_02554_ ),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_8 wire145 (.A(\soc/cpu/_01896_ ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_8 load_slew146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_6 max_cap147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_6 max_cap148 (.A(net150),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_8 load_slew149 (.A(\soc/_030_ ),
    .X(net149));
 sky130_fd_sc_hd__buf_6 max_cap150 (.A(\soc/_030_ ),
    .X(net150));
 sky130_fd_sc_hd__buf_12 load_slew151 (.A(_081_),
    .X(net151));
 sky130_fd_sc_hd__buf_16 load_slew152 (.A(\soc/cpu/cpuregs/_1677_ ),
    .X(net152));
 sky130_fd_sc_hd__buf_16 load_slew153 (.A(\soc/cpu/cpuregs/_1037_ ),
    .X(net153));
 sky130_fd_sc_hd__buf_8 max_cap154 (.A(\soc/cpu/_04116_ ),
    .X(net154));
 sky130_fd_sc_hd__buf_4 wire155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_4 load_slew156 (.A(\soc/cpu/_02705_ ),
    .X(net156));
 sky130_fd_sc_hd__buf_16 max_cap157 (.A(\soc/cpu/_02295_ ),
    .X(net157));
 sky130_fd_sc_hd__buf_16 load_slew158 (.A(\soc/cpu/_01159_ ),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_8 load_slew159 (.A(\soc/cpu/_00872_ ),
    .X(net159));
 sky130_fd_sc_hd__buf_6 max_cap160 (.A(\soc/cpu/_00872_ ),
    .X(net160));
 sky130_fd_sc_hd__buf_12 load_slew161 (.A(\soc/cpu/_00707_ ),
    .X(net161));
 sky130_fd_sc_hd__buf_12 load_slew162 (.A(\wave_gen_inst/pp ),
    .X(net162));
 sky130_fd_sc_hd__buf_16 max_cap163 (.A(\wave_gen_inst/pp ),
    .X(net163));
 sky130_fd_sc_hd__buf_6 load_slew164 (.A(net589),
    .X(net164));
 sky130_fd_sc_hd__buf_6 wire165 (.A(net588),
    .X(net165));
 sky130_fd_sc_hd__buf_2 wire166 (.A(net609),
    .X(net166));
 sky130_fd_sc_hd__buf_6 wire167 (.A(net608),
    .X(net167));
 sky130_fd_sc_hd__buf_2 wire168 (.A(net666),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 wire169 (.A(net665),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 load_slew170 (.A(net664),
    .X(net170));
 sky130_fd_sc_hd__buf_2 wire171 (.A(net663),
    .X(net171));
 sky130_fd_sc_hd__buf_2 wire172 (.A(net625),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 wire173 (.A(net624),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 wire174 (.A(net623),
    .X(net174));
 sky130_fd_sc_hd__buf_2 wire175 (.A(net633),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 wire176 (.A(net632),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 wire177 (.A(net631),
    .X(net177));
 sky130_fd_sc_hd__buf_2 wire178 (.A(net645),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 wire179 (.A(net644),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 wire180 (.A(net643),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 wire181 (.A(net572),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 wire182 (.A(net571),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 wire183 (.A(net918),
    .X(net183));
 sky130_fd_sc_hd__buf_2 wire184 (.A(net637),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 wire185 (.A(net636),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 wire186 (.A(net635),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 wire187 (.A(net586),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 wire188 (.A(net585),
    .X(net188));
 sky130_fd_sc_hd__buf_1 wire189 (.A(net584),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 wire190 (.A(net583),
    .X(net190));
 sky130_fd_sc_hd__buf_2 wire191 (.A(net641),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 wire192 (.A(net640),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 wire193 (.A(net639),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 wire194 (.A(net674),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 wire195 (.A(net673),
    .X(net195));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire196 (.A(net672),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 wire197 (.A(net671),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 wire198 (.A(net617),
    .X(net198));
 sky130_fd_sc_hd__buf_4 wire199 (.A(net616),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 wire200 (.A(net615),
    .X(net200));
 sky130_fd_sc_hd__buf_2 wire201 (.A(net670),
    .X(net201));
 sky130_fd_sc_hd__buf_2 wire202 (.A(net669),
    .X(net202));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire203 (.A(net668),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 wire204 (.A(net667),
    .X(net204));
 sky130_fd_sc_hd__buf_2 wire205 (.A(net621),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 wire206 (.A(net620),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 wire207 (.A(net619),
    .X(net207));
 sky130_fd_sc_hd__buf_2 wire208 (.A(net629),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 wire209 (.A(net628),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 wire210 (.A(net627),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 wire211 (.A(net658),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 wire212 (.A(net657),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 wire213 (.A(net656),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 wire214 (.A(net655),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 wire215 (.A(net650),
    .X(net215));
 sky130_fd_sc_hd__buf_4 wire216 (.A(net649),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 wire217 (.A(net648),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 wire218 (.A(net647),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 wire219 (.A(net581),
    .X(net219));
 sky130_fd_sc_hd__buf_4 wire220 (.A(net580),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 wire221 (.A(net920),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 wire222 (.A(net654),
    .X(net222));
 sky130_fd_sc_hd__buf_4 wire223 (.A(net653),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 wire224 (.A(net652),
    .X(net224));
 sky130_fd_sc_hd__buf_4 wire225 (.A(net651),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 wire226 (.A(net662),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 wire227 (.A(net661),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 wire228 (.A(net660),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 wire229 (.A(net659),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 wire230 (.A(net678),
    .X(net230));
 sky130_fd_sc_hd__buf_4 wire231 (.A(net677),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 wire232 (.A(net676),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 wire233 (.A(net675),
    .X(net233));
 sky130_fd_sc_hd__buf_4 wire234 (.A(net600),
    .X(net234));
 sky130_fd_sc_hd__buf_12 wire235 (.A(net916),
    .X(net235));
 sky130_fd_sc_hd__buf_4 wire236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_4 wire237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__buf_2 wire238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_1 wire239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_1 wire240 (.A(net681),
    .X(net240));
 sky130_fd_sc_hd__buf_1 wire241 (.A(net680),
    .X(net241));
 sky130_fd_sc_hd__buf_4 wire242 (.A(net679),
    .X(net242));
 sky130_fd_sc_hd__buf_4 wire243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_2 wire244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 wire245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_2 wire246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 load_slew247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_1 wire248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_1 wire249 (.A(net693),
    .X(net249));
 sky130_fd_sc_hd__buf_1 wire250 (.A(net692),
    .X(net250));
 sky130_fd_sc_hd__buf_4 wire251 (.A(net691),
    .X(net251));
 sky130_fd_sc_hd__buf_4 wire252 (.A(net606),
    .X(net252));
 sky130_fd_sc_hd__buf_12 wire253 (.A(net605),
    .X(net253));
 sky130_fd_sc_hd__buf_4 wire254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_4 wire255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__buf_2 wire256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_1 wire258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_1 wire259 (.A(net690),
    .X(net259));
 sky130_fd_sc_hd__buf_1 wire260 (.A(net689),
    .X(net260));
 sky130_fd_sc_hd__buf_4 wire261 (.A(net688),
    .X(net261));
 sky130_fd_sc_hd__buf_4 wire262 (.A(net592),
    .X(net262));
 sky130_fd_sc_hd__buf_12 wire263 (.A(net912),
    .X(net263));
 sky130_fd_sc_hd__buf_4 wire264 (.A(net603),
    .X(net264));
 sky130_fd_sc_hd__buf_16 wire265 (.A(net914),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 wire266 (.A(net613),
    .X(net266));
 sky130_fd_sc_hd__buf_12 wire267 (.A(net612),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 wire268 (.A(net611),
    .X(net268));
 sky130_fd_sc_hd__buf_4 wire269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_4 wire270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 wire271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_2 wire272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_1 wire273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_1 wire274 (.A(net687),
    .X(net274));
 sky130_fd_sc_hd__buf_4 wire275 (.A(net686),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 wire276 (.A(net685),
    .X(net276));
 sky130_fd_sc_hd__buf_4 wire277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 wire278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_8 wire279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_1 wire280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_1 wire281 (.A(net684),
    .X(net281));
 sky130_fd_sc_hd__buf_1 wire282 (.A(net683),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 wire283 (.A(net682),
    .X(net283));
 sky130_fd_sc_hd__buf_4 wire284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 wire285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 wire286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 wire287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 load_slew288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__buf_1 wire289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_1 wire290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_1 wire291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 load_slew292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_1 load_slew293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_1 wire294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_1 wire295 (.A(net700),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 wire296 (.A(net699),
    .X(net296));
 sky130_fd_sc_hd__buf_16 max_cap297 (.A(\soc/cpu/latched_stalu ),
    .X(net297));
 sky130_fd_sc_hd__buf_16 load_slew298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_12 load_slew299 (.A(net301),
    .X(net299));
 sky130_fd_sc_hd__buf_12 load_slew300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_16 load_slew301 (.A(\soc/cpu/cpuregs_raddr2[4] ),
    .X(net301));
 sky130_fd_sc_hd__buf_16 load_slew302 (.A(net304),
    .X(net302));
 sky130_fd_sc_hd__buf_16 max_cap303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_16 load_slew304 (.A(\soc/cpu/cpuregs_raddr2[3] ),
    .X(net304));
 sky130_fd_sc_hd__buf_12 load_slew305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_16 load_slew306 (.A(net309),
    .X(net306));
 sky130_fd_sc_hd__buf_16 wire307 (.A(net309),
    .X(net307));
 sky130_fd_sc_hd__buf_16 load_slew308 (.A(net310),
    .X(net308));
 sky130_fd_sc_hd__buf_16 max_cap309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_16 load_slew310 (.A(\soc/cpu/cpuregs_raddr2[2] ),
    .X(net310));
 sky130_fd_sc_hd__buf_16 load_slew311 (.A(\soc/cpu/cpuregs_raddr2[2] ),
    .X(net311));
 sky130_fd_sc_hd__buf_16 load_slew312 (.A(\soc/cpu/cpuregs_raddr2[2] ),
    .X(net312));
 sky130_fd_sc_hd__buf_16 wire313 (.A(net315),
    .X(net313));
 sky130_fd_sc_hd__buf_16 wire314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_16 wire315 (.A(\soc/cpu/cpuregs_raddr2[1] ),
    .X(net315));
 sky130_fd_sc_hd__buf_16 max_cap316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_16 load_slew317 (.A(net320),
    .X(net317));
 sky130_fd_sc_hd__buf_12 load_slew318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_16 load_slew319 (.A(net324),
    .X(net319));
 sky130_fd_sc_hd__buf_16 load_slew320 (.A(net324),
    .X(net320));
 sky130_fd_sc_hd__buf_16 max_cap321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__buf_16 wire322 (.A(net324),
    .X(net322));
 sky130_fd_sc_hd__buf_12 load_slew323 (.A(net326),
    .X(net323));
 sky130_fd_sc_hd__buf_16 load_slew324 (.A(net326),
    .X(net324));
 sky130_fd_sc_hd__buf_16 wire325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__buf_16 load_slew326 (.A(\soc/cpu/cpuregs_raddr2[0] ),
    .X(net326));
 sky130_fd_sc_hd__buf_16 load_slew327 (.A(net329),
    .X(net327));
 sky130_fd_sc_hd__buf_16 wire328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_16 wire329 (.A(\soc/cpu/cpuregs_raddr1[4] ),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_16 load_slew330 (.A(net332),
    .X(net330));
 sky130_fd_sc_hd__buf_16 load_slew331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__buf_16 load_slew332 (.A(\soc/cpu/cpuregs_raddr1[3] ),
    .X(net332));
 sky130_fd_sc_hd__buf_16 load_slew333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_16 load_slew334 (.A(\soc/cpu/cpuregs_raddr1[2] ),
    .X(net334));
 sky130_fd_sc_hd__buf_12 load_slew335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__buf_16 load_slew336 (.A(\soc/cpu/cpuregs_raddr1[2] ),
    .X(net336));
 sky130_fd_sc_hd__buf_16 load_slew337 (.A(net340),
    .X(net337));
 sky130_fd_sc_hd__buf_16 load_slew338 (.A(net340),
    .X(net338));
 sky130_fd_sc_hd__buf_16 max_cap339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__buf_16 load_slew340 (.A(\soc/cpu/cpuregs_raddr1[2] ),
    .X(net340));
 sky130_fd_sc_hd__buf_12 load_slew341 (.A(net343),
    .X(net341));
 sky130_fd_sc_hd__buf_16 load_slew342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__buf_16 wire343 (.A(\soc/cpu/cpuregs_raddr1[1] ),
    .X(net343));
 sky130_fd_sc_hd__buf_16 load_slew344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_16 load_slew345 (.A(net348),
    .X(net345));
 sky130_fd_sc_hd__buf_16 max_cap346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_16 load_slew347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_16 load_slew348 (.A(net353),
    .X(net348));
 sky130_fd_sc_hd__buf_16 wire349 (.A(net353),
    .X(net349));
 sky130_fd_sc_hd__buf_12 load_slew350 (.A(net352),
    .X(net350));
 sky130_fd_sc_hd__buf_16 max_cap351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_16 load_slew352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__buf_16 wire353 (.A(\soc/cpu/cpuregs_raddr1[0] ),
    .X(net353));
 sky130_fd_sc_hd__buf_2 wire354 (.A(net524),
    .X(net354));
 sky130_fd_sc_hd__buf_2 wire355 (.A(net523),
    .X(net355));
 sky130_fd_sc_hd__buf_1 wire356 (.A(net522),
    .X(net356));
 sky130_fd_sc_hd__buf_2 wire357 (.A(net521),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_4 wire358 (.A(net520),
    .X(net358));
 sky130_fd_sc_hd__buf_2 wire359 (.A(net518),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 wire360 (.A(net517),
    .X(net360));
 sky130_fd_sc_hd__buf_1 wire361 (.A(net516),
    .X(net361));
 sky130_fd_sc_hd__buf_2 wire362 (.A(net515),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 wire363 (.A(net514),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 wire364 (.A(net902),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_8 wire365 (.A(net900),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 wire366 (.A(net508),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 wire367 (.A(net507),
    .X(net367));
 sky130_fd_sc_hd__buf_1 wire368 (.A(net506),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 load_slew369 (.A(net505),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 wire370 (.A(net504),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 wire371 (.A(net502),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 wire372 (.A(net501),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 wire373 (.A(net500),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_4 wire374 (.A(net721),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 wire375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 wire376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_1 wire377 (.A(net598),
    .X(net377));
 sky130_fd_sc_hd__buf_1 wire378 (.A(net597),
    .X(net378));
 sky130_fd_sc_hd__buf_1 wire379 (.A(net596),
    .X(net379));
 sky130_fd_sc_hd__buf_1 wire380 (.A(net595),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_4 wire381 (.A(net594),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 wire382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 wire383 (.A(net531),
    .X(net383));
 sky130_fd_sc_hd__buf_1 wire384 (.A(net530),
    .X(net384));
 sky130_fd_sc_hd__buf_1 wire385 (.A(net529),
    .X(net385));
 sky130_fd_sc_hd__buf_1 wire386 (.A(net528),
    .X(net386));
 sky130_fd_sc_hd__buf_2 wire387 (.A(net527),
    .X(net387));
 sky130_fd_sc_hd__buf_4 wire388 (.A(net526),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 wire389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 wire390 (.A(net537),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 wire391 (.A(net536),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 load_slew392 (.A(net535),
    .X(net392));
 sky130_fd_sc_hd__buf_1 wire393 (.A(net534),
    .X(net393));
 sky130_fd_sc_hd__buf_2 wire394 (.A(net533),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_4 wire395 (.A(net532),
    .X(net395));
 sky130_fd_sc_hd__buf_12 load_slew396 (.A(\soc/cpu/irq_state[0] ),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 wire397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 wire398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_1 wire399 (.A(net545),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_8 wire400 (.A(net558),
    .X(net400));
 sky130_fd_sc_hd__buf_2 wire401 (.A(net577),
    .X(net401));
 sky130_fd_sc_hd__buf_4 wire402 (.A(net576),
    .X(net402));
 sky130_fd_sc_hd__buf_2 wire403 (.A(net575),
    .X(net403));
 sky130_fd_sc_hd__buf_1 wire404 (.A(net574),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_4 wire405 (.A(net563),
    .X(net405));
 sky130_fd_sc_hd__buf_4 wire406 (.A(net562),
    .X(net406));
 sky130_fd_sc_hd__buf_2 wire407 (.A(net561),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 wire408 (.A(net560),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_4 wire409 (.A(net568),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 wire410 (.A(net567),
    .X(net410));
 sky130_fd_sc_hd__buf_2 wire411 (.A(net566),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 wire412 (.A(net565),
    .X(net412));
 sky130_fd_sc_hd__buf_16 load_slew413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__buf_12 load_slew414 (.A(net801),
    .X(net414));
 sky130_fd_sc_hd__buf_16 wire415 (.A(\soc/ram_ready ),
    .X(net415));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06662__416  (.LO(net416));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06664__417  (.LO(net417));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06666__418  (.LO(net418));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06657__420  (.LO(net420));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06659__421  (.LO(net421));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06668__422  (.LO(net422));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06670__423  (.LO(net423));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06672__424  (.LO(net424));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06675__425  (.LO(net425));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06677__426  (.LO(net426));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06679__427  (.LO(net427));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06681__428  (.LO(net428));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06684__429  (.LO(net429));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06686__430  (.LO(net430));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06688__431  (.LO(net431));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06690__432  (.LO(net432));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06692__433  (.LO(net433));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06694__434  (.LO(net434));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06697__435  (.LO(net435));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06699__436  (.LO(net436));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06701__437  (.LO(net437));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06703__438  (.LO(net438));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06706__439  (.LO(net439));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06708__440  (.LO(net440));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06710__441  (.LO(net441));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06712__442  (.LO(net442));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06714__443  (.LO(net443));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06716__444  (.LO(net444));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_06718__445  (.LO(net445));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_05182__446  (.LO(net446));
 sky130_fd_sc_hd__conb_1 \soc/cpu/_05231__447  (.LO(net447));
 sky130_fd_sc_hd__conb_1 \soc/_243__449  (.LO(net449));
 sky130_fd_sc_hd__conb_1 \soc/_252__450  (.LO(net450));
 sky130_fd_sc_hd__conb_1 \soc/_252__451  (.LO(net451));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/_0564__452  (.LO(net452));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/_0565__453  (.LO(net453));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/_0759__454  (.LO(net454));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/_0764__455  (.LO(net455));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/_0962__456  (.LO(net456));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/_0971__457  (.LO(net457));
 sky130_fd_sc_hd__conb_1 \soc/_332__459  (.LO(net459));
 sky130_fd_sc_hd__conb_1 \soc/_369__460  (.LO(net460));
 sky130_fd_sc_hd__conb_1 \soc/_375__461  (.LO(net461));
 sky130_fd_sc_hd__conb_1 \soc/_381__462  (.LO(net462));
 sky130_fd_sc_hd__conb_1 \soc/_389__463  (.LO(net463));
 sky130_fd_sc_hd__conb_1 \soc/_444__464  (.LO(net464));
 sky130_fd_sc_hd__conb_1 \soc/_450__465  (.LO(net465));
 sky130_fd_sc_hd__conb_1 \soc/_456__466  (.LO(net466));
 sky130_fd_sc_hd__conb_1 \soc/_462__467  (.LO(net467));
 sky130_fd_sc_hd__conb_1 \soc/_468__468  (.LO(net468));
 sky130_fd_sc_hd__conb_1 \soc/_474__469  (.LO(net469));
 sky130_fd_sc_hd__conb_1 \soc/_480__470  (.LO(net470));
 sky130_fd_sc_hd__conb_1 \soc/_486__471  (.LO(net471));
 sky130_fd_sc_hd__conb_1 \soc/spimemio/xfer/_364__472  (.LO(net472));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3056__475  (.HI(net475));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3089__476  (.HI(net476));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3120__477  (.HI(net477));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3144__478  (.HI(net478));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3205__479  (.HI(net479));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3231__480  (.HI(net480));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3250__481  (.HI(net481));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3272__482  (.HI(net482));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3273__483  (.HI(net483));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3308__484  (.HI(net484));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3347__485  (.HI(net485));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3375__486  (.HI(net486));
 sky130_fd_sc_hd__conb_1 \wave_gen_inst/_3377__487  (.HI(net487));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0743__489  (.A(clknet_leaf_73_clk),
    .Y(net489));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0743__490  (.A(clknet_leaf_73_clk),
    .Y(net490));
 sky130_fd_sc_hd__inv_1 \soc/spimemio/_0743__491  (.A(clknet_leaf_73_clk),
    .Y(net491));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_1_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_2_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_3_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_4_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_5_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_6_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_7_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_8_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_9_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_10_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_11_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_12_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_13_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_14_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_15_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_16_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_17_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_18_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_19_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_20_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_21_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_22_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_23_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_24_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_25_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_26_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_27_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_28_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_29_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_30_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_31_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_32_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_33_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_34_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_35_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_36_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_37_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_38_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_39_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_40_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_41_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_42_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_43_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_44_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_45_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_46_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_47_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_48_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_49_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_50_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_51_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_52_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_53_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_54_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_55_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_56_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_57_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_58_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_59_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_60_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_61_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_62_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_63_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_65_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_66_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_67_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_68_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_69_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_70_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_71_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_72_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_73_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_74_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_75_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_76_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_77_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_78_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_79_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_80_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_81_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_82_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_83_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_84_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_85_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_86_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_87_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_88_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_89_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_90_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_91_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_92_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_93_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_leaf_94_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\iomem_addr[25] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(net766),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(net909),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(net67),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net899),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(net901),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net364),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net720),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net374),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(net373),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(net372),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(net371),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(net938),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net370),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(net369),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(net368),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(net367),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(net366),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\soc/simpleuart/recv_divcnt[19] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net539),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(net922),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\soc/simpleuart/_0112_ ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(net940),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(net363),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net362),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net361),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(net360),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net359),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net945),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(net358),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net357),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(net356),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(net355),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(net354),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\iomem_addr[3] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(net388),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net387),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net386),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(net385),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net384),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\iomem_addr[2] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(net395),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net394),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(net393),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(net392),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net391),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\soc/simpleuart/recv_divcnt[18] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\soc/simpleuart/_0641_ ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(net511),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\soc/simpleuart/_0646_ ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\soc/simpleuart/_0648_ ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\soc/simpleuart/_0113_ ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(net557),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(net559),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\soc/_011_ ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\soc/simpleuart/_0335_ ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\soc/simpleuart/_0000_ ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\soc/simpleuart/recv_divcnt[17] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\soc/simpleuart/_0439_ ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\soc/simpleuart/_0448_ ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\soc/simpleuart/_0472_ ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\soc/simpleuart/_0485_ ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\soc/simpleuart/_0567_ ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\soc/simpleuart/_0607_ ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\soc/simpleuart/_0114_ ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\iomem_wstrb[3] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(net544),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net400),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(net934),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(net408),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(net407),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(net406),
    .X(net563));
 sky130_fd_sc_hd__buf_2 hold564 (.A(net405),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(net937),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(net412),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(net411),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(net410),
    .X(net568));
 sky130_fd_sc_hd__buf_2 hold569 (.A(net409),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(net917),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(net183),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(net182),
    .X(net572));
 sky130_fd_sc_hd__buf_2 hold573 (.A(net181),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net936),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(net404),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(net403),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(net402),
    .X(net577));
 sky130_fd_sc_hd__buf_2 hold578 (.A(net401),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(net919),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(net221),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(net220),
    .X(net581));
 sky130_fd_sc_hd__buf_2 hold582 (.A(net219),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net935),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(net190),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(net189),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(net188),
    .X(net586));
 sky130_fd_sc_hd__buf_2 hold587 (.A(net187),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(net924),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(net165),
    .X(net589));
 sky130_fd_sc_hd__buf_2 hold590 (.A(net164),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net911),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(net263),
    .X(net592));
 sky130_fd_sc_hd__buf_2 hold593 (.A(net262),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\iomem_addr[4] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(net381),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(net380),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net379),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(net378),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(net915),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(net235),
    .X(net600));
 sky130_fd_sc_hd__buf_2 hold601 (.A(net234),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(net913),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(net265),
    .X(net603));
 sky130_fd_sc_hd__buf_2 hold604 (.A(net264),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(net782),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net253),
    .X(net606));
 sky130_fd_sc_hd__buf_2 hold607 (.A(net252),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(net926),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(net167),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 hold610 (.A(net166),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(net932),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(net268),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(net267),
    .X(net613));
 sky130_fd_sc_hd__buf_2 hold614 (.A(net266),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(net930),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(net200),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(net199),
    .X(net617));
 sky130_fd_sc_hd__buf_2 hold618 (.A(net198),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(net929),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(net207),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(net206),
    .X(net621));
 sky130_fd_sc_hd__buf_2 hold622 (.A(net205),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(net928),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(net174),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(net173),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_4 hold626 (.A(net172),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(net931),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(net210),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(net209),
    .X(net629));
 sky130_fd_sc_hd__buf_2 hold630 (.A(net208),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(net823),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(net177),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(net176),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_4 hold634 (.A(net175),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(net815),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net186),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(net185),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_4 hold638 (.A(net184),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(net806),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(net193),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(net192),
    .X(net641));
 sky130_fd_sc_hd__buf_2 hold642 (.A(net191),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(net933),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(net180),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(net179),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_4 hold646 (.A(net178),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\iomem_wdata[15] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(net218),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(net217),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(net216),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\iomem_wdata[13] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(net225),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(net224),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(net223),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\iomem_wdata[16] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(net214),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(net213),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(net212),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\iomem_wdata[12] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(net229),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net228),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(net227),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\iomem_wdata[29] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net171),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(net170),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(net169),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\iomem_wdata[19] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(net204),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(net203),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(net202),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\iomem_wdata[21] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(net197),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(net196),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(net195),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\iomem_wdata[11] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(net233),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(net232),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(net231),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\iomem_wdata[9] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(net242),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(net241),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\iomem_wdata[1] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(net283),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(net282),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\iomem_wdata[2] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(net276),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net275),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\iomem_wdata[6] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(net261),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(net260),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\iomem_wdata[8] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(net251),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(net250),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\iomem_addr[23] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\soc/spimemio/_0366_ ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\soc/spimemio/_0048_ ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(net949),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\soc/cpu/_02847_ ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\iomem_wdata[0] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(net296),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\iomem_addr[27] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_084_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_182_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\gpio[30] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_123_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_044_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(net723),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\iomem_addr[14] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\soc/spimemio/_0480_ ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\soc/spimemio/buffer[11] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\soc/spimemio/_0396_ ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\soc/spimemio/_0068_ ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\iomem_addr[15] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\iomem_addr[10] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\soc/spimemio/_0338_ ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\soc/spimemio/_0035_ ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\iomem_addr[30] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_079_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_126_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\iomem_addr[5] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(net499),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\soc/spimemio/dout_tag[2] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\soc/simpleuart/recv_divcnt[20] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\iomem_addr[18] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\soc/_013_ ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\soc/_017_ ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\soc/_001_ ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\soc/spimemio/rd_addr[16] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\soc/spimemio/_0210_ ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\soc/spimemio/_0238_ ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\soc/spimemio/_0239_ ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\soc/spimemio/_0240_ ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\soc/spimemio/_0244_ ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\soc/spimemio/_0009_ ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\soc/spimemio/softreset ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\iomem_addr[16] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\soc/spimemio/_0448_ ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\soc/spimemio/_0091_ ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\iomem_addr[29] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\soc/_018_ ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\soc/_021_ ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\soc/_037_ ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(net135),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\iomem_addr[11] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\soc/spimemio/_0036_ ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\soc/spimemio/config_cont ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\soc/spimemio/rd_addr[2] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\soc/spimemio/_0218_ ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\soc/spimemio/_0030_ ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\soc/spimemio/rd_addr[3] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\soc/cpu/instr_sltiu ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\soc/cpu/_00035_ ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\soc/spimemio/dout_data[1] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\soc/cpu/pcpi_rs2 [22]),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\soc/cpu/_01997_ ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\soc/spimemio_cfgreg_do[19] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(net37),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_091_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_016_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\soc/cpu/count_instr[13] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\soc/cpu/_04619_ ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\soc/cpu/_00420_ ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\iomem_addr[31] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\soc/_019_ ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\soc/_040_ ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\soc/_041_ ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(net493),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net26),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(_090_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_015_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\iomem_addr[12] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\soc/simpleuart/send_dummy ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\soc/cpu/mem_la_wdata [7]),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\soc/cpu/_01829_ ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\soc/cpu/alu_out[7] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\soc/cpu/mem_la_wdata [6]),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\soc/cpu/pcpi_rs2 [11]),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\soc/cpu/cpu_state[0] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\iomem_addr[17] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\soc/cpu/pcpi_rs2 [8]),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\soc/cpu/pcpi_rs2 [9]),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(net927),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\soc/spimemio/rd_addr[6] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\soc/cpu/decoder_pseudo_trigger ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\soc/cpu/count_instr[12] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\soc/cpu/_04616_ ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\iomem_rdata[27] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\soc/cpu/mem_la_wdata [6]),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\soc/cpu/count_cycle[43] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\soc/cpu/_04077_ ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\soc/cpu/_00324_ ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\soc/cpu/count_instr[43] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\soc/cpu/_04716_ ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\soc/cpu/_00458_ ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\soc/cpu/count_cycle[42] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(net43),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_095_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\soc/cpu/count_instr[11] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\soc/cpu/mem_do_prefetch ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\soc/cpu/_00842_ ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\soc/cpu/cpu_state[2] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\soc/cpu/instr_sltu ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\wave_gen_inst/param1[4] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\soc/cpu/reg_sh[0] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\iomem_rdata[21] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\iomem_wdata[22] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\soc/cpu/cpu_state[2] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(iomem_ready),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\iomem_addr[26] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_098_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\soc/cpu/count_instr[42] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\soc/cpu/_04692_ ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\wave_gen_inst/counter[19] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\wave_gen_inst/counter[21] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\iomem_wdata[24] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\iomem_rdata[29] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\wave_gen_inst/counter[22] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\wave_gen_inst/counter[25] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\soc/cpu/cpu_state[1] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\soc/cpu/_00401_ ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\wave_gen_inst/param1[1] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\soc/spimemio/rd_valid ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\iomem_wdata[27] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\soc/spimemio/rd_addr[13] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\soc/spimemio/_0140_ ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\soc/spimemio/_0146_ ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\soc/spimemio/_0147_ ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\soc/spimem_ready ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\wave_gen_inst/counter[9] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\wave_gen_inst/_1078_ ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\wave_gen_inst/_1087_ ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\wave_gen_inst/_1092_ ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\iomem_rdata[28] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\soc/cpu/reg_pc[8] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\soc/cpu/pcpi_rs1 [7]),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\soc/cpu/_00188_ ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\reset_cnt[3] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_078_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\wave_gen_inst/param1[3] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\soc/cpu/reg_pc[8] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\soc/spimemio/buffer[20] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(net925),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\wave_gen_inst/counter[1] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\wave_gen_inst/_0920_ ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\wave_gen_inst/_1507_ ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\wave_gen_inst/counter[10] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\wave_gen_inst/_1103_ ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\soc/cpu/mem_la_wdata [1]),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\wave_gen_inst/param1[2] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\soc/cpu/is_alu_reg_reg ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\soc/cpu/pcpi_rs1 [1]),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\soc/cpu/mem_rdata_q[14] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\soc/cpu/decoded_imm[29] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\soc/cpu/decoded_imm[28] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\soc/cpu/mem_la_wdata [2]),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\soc/cpu/irq_pending[2] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\soc/cpu/decoded_imm[3] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\iomem_rdata[17] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\iomem_rdata[22] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\soc/cpu/pcpi_rs1 [5]),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\soc/cpu/reg_out[0] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\soc/cpu/reg_next_pc[5] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\soc/spimemio/din_qspi ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\soc/spimemio/rd_addr[22] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\soc/spimemio/_0189_ ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\soc/cpu/irq_mask[18] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(net923),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\iomem_rdata[26] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\gpio[24] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\soc/spimemio/xfer/xfer_tag[3] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\soc/spimemio/xfer/xfer_tag[2] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\soc/cpu/decoded_imm[10] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\soc/cpu/reg_pc[4] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\soc/cpu/decoded_imm[9] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\soc/cpu/mem_rdata_q[27] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\soc/cpu/irq_mask[0] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\soc/cpu/_00001_ ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\soc/cpu/decoded_imm[31] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\soc/cpu/decoded_imm[12] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\wave_gen_inst/counter[7] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\soc/cpu/pcpi_rs1 [19]),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\wave_gen_inst/counter[24] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\soc/cpu/latched_compr ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\soc/spimemio/rd_addr[18] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\soc/cpu/timer[0] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\soc/spimemio/dout_data[4] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\soc/cpu/irq_mask[11] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\soc/cpu/pcpi_rs1 [17]),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\soc/cpu/decoded_imm[20] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\soc/cpu/decoded_imm[19] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\soc/spimemio/xfer/xfer_tag[1] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\soc/cpu/mem_state[0] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\soc/cpu/pcpi_rs1 [21]),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\soc/spimemio/xfer/xfer_tag[0] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\soc/cpu/pcpi_rs1 [23]),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\iomem_rdata[31] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\soc/cpu/pcpi_rs1 [25]),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\soc/cpu/decoded_rd[4] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\iomem_addr[7] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(net496),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(net365),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(net497),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\soc/mem_valid ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\soc/_033_ ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\soc/_034_ ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net137),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\soc/_039_ ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\soc/mem_ready ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\soc/_003_ ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(net494),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\iomem_wdata[5] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(net591),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\iomem_wdata[4] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(net602),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\iomem_wdata[10] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(net599),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\iomem_wdata[25] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(net570),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\iomem_wdata[14] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(net579),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\soc/simpleuart/recv_divcnt[21] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\soc/simpleuart/_0647_ ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\iomem_wdata[31] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(net867),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\iomem_wdata[30] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(net842),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\iomem_wdata[7] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\iomem_wdata[28] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\iomem_wdata[18] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\iomem_wdata[20] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\iomem_wdata[17] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\iomem_wdata[3] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\iomem_wdata[26] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\iomem_wstrb[1] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\iomem_wdata[23] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\iomem_wstrb[2] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\iomem_wstrb[0] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\iomem_addr[6] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\soc/spimemio/rd_addr[21] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\iomem_addr[8] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\iomem_addr[26] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_163_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\wave_gen_inst/counter[10] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\reset_cnt[1] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\iomem_addr[9] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\iomem_addr[17] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\iomem_addr[14] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\soc/cpu/decoded_imm[12] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\soc/cpu/is_alu_reg_imm ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\soc/cpu/mem_rdata_q[14] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\soc/cpu/mem_rdata_q[13] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\soc/cpu/is_sb_sh_sw ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\soc/cpu/is_lb_lh_lw_lbu_lhu ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\soc/cpu/is_beq_bne_blt_bge_bltu_bgeu ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\soc/cpu/cpu_state[2] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\soc/cpu/mem_rdata_q[13] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\soc/cpu/mem_rdata_q[24] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\iomem_rdata[19] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\wave_gen_inst/counter[9] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\soc/cpu/irq_pending[6] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\soc/cpu/_03540_ ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\soc/cpu/cpuregs_raddr2[4] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\soc/cpu/cpuregs_raddr2[3] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\soc/cpu/decoded_imm_j[6] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\soc/cpu/_02786_ ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\iomem_rdata[25] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\soc/cpu/pcpi_rs1 [3]),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\wave_gen_inst/counter[10] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\soc/cpu/mem_la_wdata [1]),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\soc/spimemio/dout_data[2] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\soc/spimemio/dout_data[4] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\soc/cpu/pcpi_rs2 [22]),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\wave_gen_inst/param1[4] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\soc/cpu/count_instr[41] ),
    .X(net974));
endmodule
